module LSHIFT2(input [15:0] entrada, output [17:0] saida);
	assign saida = entrada << 2;
endmodule