.include transmissiongate2.spi

x1 10 11 20 30 40 transmissiongate2

v1 10 30 sine(0.9 0.9 2G 0 0 0)
v3 20 30 1.8V
v5 30 0 0V DC
v6 11 30 pulse(0 1.8 0ns 1ps 1ps 2ns 4ns)

r1 40 30 100k

.tran 1ps 8000ps

.model tp pmos level=54
.model tn nmos level=54

.end
