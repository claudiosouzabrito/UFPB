* Spice description of inversores
* Spice driver version 507442696
* Date ( dd/mm/yyyy hh:mm:ss ):  3/07/2019 at 23:35:57

* INTERF a vdd vss y y1 y2 


.subckt inversores 9 30 70 53 37 2 
* NET 2 = y2
* NET 9 = a
* NET 30 = vdd
* NET 37 = y1
* NET 53 = y
* NET 70 = vss
Mtr_00006 21 43 4 30 tp L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00005 20 59 42 30 tp L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00004 19 14 58 30 tp L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_00003 1 36 73 70 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00002 33 52 69 70 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00001 49 11 65 70 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
R6_1 1 3 0.001
R6_2 4 5 0.001
R6_3 5 6 0.1
C6_31 5 70 3.5e-16
C6_32 6 70 3.5e-16
R6_4 2 5 0.8
C6_41 2 70 2.38e-15
C6_42 5 70 2.38e-15
R6_5 3 2 0.4
C6_51 3 70 1.26e-15
C6_52 2 70 1.26e-15
R5_1 13 12 0.001
R5_2 12 16 0.7
C5_21 12 70 2.17e-15
C5_22 16 70 2.17e-15
R5_3 9 12 0.3
C5_31 9 70 8.4e-16
C5_32 12 70 8.4e-16
R5_4 10 9 0.3
C5_41 10 70 1.05e-15
C5_42 9 70 1.05e-15
R5_5 13 15 200
C5_51 13 70 6e-16
C5_52 15 70 6e-16
R5_6 15 14 450
C5_61 15 70 1.425e-15
C5_62 14 70 1.425e-15
R5_7 11 15 550
C5_71 11 70 1.65e-15
C5_72 15 70 1.65e-15
R4_1 19 22 0.001
R4_2 21 27 0.001
R4_3 20 26 0.001
R4_4 28 29 0.001
C4_41 28 70 8.4e-16
C4_42 29 70 8.4e-16
R4_5 27 28 0.1
C4_51 27 70 1.44e-15
C4_52 28 70 1.44e-15
R4_6 25 27 0.1
C4_61 25 70 2.64e-15
C4_62 27 70 2.64e-15
R4_7 25 30 0.001
C4_71 25 70 7.2e-16
C4_72 30 70 7.2e-16
R4_8 26 30 0.001
C4_81 26 70 7.2e-16
C4_82 30 70 7.2e-16
R4_9 23 26 0.1
C4_91 23 70 2.64e-15
C4_92 26 70 2.64e-15
R4_10 22 23 0.1
C4_101 22 70 1.44e-15
C4_102 23 70 1.44e-15
R4_11 24 22 0.001
C4_111 24 70 6e-16
C4_112 22 70 6e-16
R3_1 33 34 0.001
R3_2 42 44 0.001
R3_3 40 39 0.001
R3_4 41 43 450
C3_41 41 70 1.425e-15
C3_42 43 70 1.425e-15
R3_5 36 41 550
C3_51 36 70 1.65e-15
C3_52 41 70 1.65e-15
R3_6 40 41 200
C3_61 40 70 6e-16
C3_62 41 70 6e-16
R3_7 39 46 0.7
C3_71 39 70 2.17e-15
C3_72 46 70 2.17e-15
R3_8 35 39 0.6
C3_81 35 70 1.89e-15
C3_82 39 70 1.89e-15
R3_9 38 39 1
C3_91 38 70 1.2075e-15
C3_92 39 70 1.2075e-15
R3_10 44 45 0.1
C3_101 44 70 3.5e-16
C3_102 45 70 3.5e-16
R3_11 38 44 0.6
C3_111 38 70 1.82e-15
C3_112 44 70 1.82e-15
R3_12 37 38 0.2
C3_121 37 70 5.6e-16
C3_122 38 70 5.6e-16
R3_13 34 37 0.4
C3_131 34 70 1.26e-15
C3_132 37 70 1.26e-15
R2_1 49 50 0.001
R2_2 58 60 0.001
R2_3 56 55 0.001
R2_4 57 59 450
C2_41 57 70 1.425e-15
C2_42 59 70 1.425e-15
R2_5 52 57 550
C2_51 52 70 1.65e-15
C2_52 57 70 1.65e-15
R2_6 56 57 200
C2_61 56 70 6e-16
C2_62 57 70 6e-16
R2_7 55 62 0.7
C2_71 55 70 2.17e-15
C2_72 62 70 2.17e-15
R2_8 51 55 0.6
C2_81 51 70 1.89e-15
C2_82 55 70 1.89e-15
R2_9 54 55 1
C2_91 54 70 1.2075e-15
C2_92 55 70 1.2075e-15
R2_10 60 61 0.1
C2_101 60 70 3.5e-16
C2_102 61 70 3.5e-16
R2_11 54 60 0.6
C2_111 54 70 1.82e-15
C2_112 60 70 1.82e-15
R2_12 53 54 0.2
C2_121 53 70 5.6e-16
C2_122 54 70 5.6e-16
R2_13 50 53 0.4
C2_131 50 70 1.26e-15
C2_132 53 70 1.26e-15
R1_1 69 71 0.001
R1_2 73 74 0.001
R1_3 65 67 0.001
R1_4 75 76 0.001
C1_41 75 70 8.4e-16
C1_42 76 70 8.4e-16
R1_5 74 75 0.1
C1_51 74 70 1.44e-15
C1_52 75 70 1.44e-15
R1_6 72 74 0.1
C1_61 72 70 2.64e-15
C1_62 74 70 2.64e-15
R1_7 72 70 0.001
C1_71 72 70 7.2e-16
C1_72 70 70 7.2e-16
R1_8 71 70 0.001
C1_81 71 70 7.2e-16
C1_82 70 70 7.2e-16
R1_9 66 71 0.1
C1_91 66 70 2.4e-15
C1_92 71 70 2.4e-15
R1_10 67 66 0.1
C1_101 67 70 1.68e-15
C1_102 66 70 1.68e-15
R1_11 68 67 0.001
C1_111 68 70 6e-16
C1_112 67 70 6e-16
.ends inversores

