* Spice description of transmissiongate
* Spice driver version 1891989000
* Date ( dd/mm/yyyy hh:mm:ss ): 26/08/2019 at 21:36:37

* INTERF a s vdd vss y1 y2 


.subckt transmissiongate 5 1 2 7 3 4 
* NET 1 = s
* NET 2 = vdd
* NET 3 = y1
* NET 4 = y2
* NET 5 = a
* NET 6 = inversor_1.nq
* NET 7 = vss
Mtr_00006 6 1 2 2 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00005 2 1 6 2 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00004 5 1 3 2 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00003 7 1 6 7 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00002 7 1 6 7 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00001 5 6 4 7 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
C7 1 7 3.776e-14
C6 2 7 1.015e-14
C5 3 7 1.94e-15
C4 4 7 1.94e-15
C3 5 7 7.33e-15
C2 6 7 3.092e-14
C1 7 7 9.59e-15
.ends transmissiongate

