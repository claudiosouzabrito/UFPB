* Spice description of 2faseclk
* Spice driver version 973764104
* Date ( dd/mm/yyyy hh:mm:ss ): 19/08/2019 at 13:53:21

* INTERF clk q qb vdd vss vss 


.subckt 2faseclk 85 48 115 137 193 209 
* NET 4 = inv3.nq
* NET 21 = nand2.nq
* NET 48 = q
* NET 63 = inv2.nq
* NET 85 = clk
* NET 115 = qb
* NET 137 = vdd
* NET 154 = nand1.nq
* NET 171 = inv1.nq
* NET 193 = vss
* NET 209 = vss
Mtr_00018 175 84 127 137 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00017 162 176 128 137 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00016 129 106 162 137 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00015 70 161 130 137 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00014 40 69 131 137 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00013 116 11 151 137 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00012 4 25 150 137 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00011 21 54 148 137 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00010 149 88 21 137 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00009 189 80 171 193 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00008 192 174 186 193 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00007 186 102 154 193 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00006 197 157 63 193 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00005 201 66 38 193 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00004 215 15 123 193 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00003 211 32 16 193 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00002 206 59 1 193 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00001 1 96 31 193 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
R11_1 4 5 0.001
R11_2 4 12 0.001
R11_3 5 6 0.001
R11_4 16 17 0.001
R11_5 9 8 0.001
R11_6 14 13 0.001
R11_7 14 15 500
C11_71 14 193 1.5e-15
C11_72 15 193 1.5e-15
R11_8 11 14 600
C11_81 11 193 1.875e-15
C11_82 14 193 1.875e-15
R11_9 13 18 0.5
C11_91 13 193 1.47e-15
C11_92 18 193 1.47e-15
R11_10 8 13 0.7
C11_101 8 193 2.1e-15
C11_102 13 193 2.1e-15
R11_11 10 8 0.2
C11_111 10 193 7.7e-16
C11_112 8 193 7.7e-16
R11_12 6 9 0.25
C11_121 6 193 1.2e-15
C11_122 9 193 1.2e-15
R11_13 12 17 1
C11_131 12 193 2.8e-15
C11_132 17 193 2.8e-15
R11_14 5 12 0.2
C11_141 5 193 7e-16
C11_142 12 193 7e-16
R11_15 7 5 0.2
C11_151 7 193 7.7e-16
C11_152 5 193 7.7e-16
R10_1 21 22 0.001
R10_2 21 23 0.001
R10_3 22 24 0.001
R10_4 31 34 0.001
R10_5 27 26 0.001
R10_6 29 30 0.001
R10_7 29 32 500
C10_71 29 193 1.5e-15
C10_72 32 193 1.5e-15
R10_8 25 29 600
C10_81 25 193 1.875e-15
C10_82 29 193 1.875e-15
R10_9 30 35 0.5
C10_91 30 193 1.47e-15
C10_92 35 193 1.47e-15
R10_10 26 30 0.7
C10_101 26 193 2.1e-15
C10_102 30 193 2.1e-15
R10_11 28 26 0.2
C10_111 28 193 7.7e-16
C10_112 26 193 7.7e-16
R10_12 24 27 0.35
C10_121 24 193 1.8e-15
C10_122 27 193 1.8e-15
R10_13 33 34 0.2
C10_131 33 193 5.6e-16
C10_132 34 193 5.6e-16
R10_14 22 33 1.2
C10_141 22 193 3.5e-15
C10_142 33 193 3.5e-15
R10_15 23 22 0.2
C10_151 23 193 7e-16
C10_152 22 193 7e-16
R9_1 38 39 0.001
R9_2 40 41 0.001
R9_3 49 48 0.001
R9_4 40 42 0.001
R9_5 49 50 0.001
R9_6 52 51 0.001
R9_7 44 43 0.001
R9_8 56 55 0.001
R9_9 55 57 0.001
R9_10 54 58 0.001
R9_11 54 59 1150
C9_111 54 193 3.5625e-15
C9_112 59 193 3.5625e-15
R9_12 58 60 1
C9_121 58 193 2.87e-15
C9_122 60 193 2.87e-15
R9_13 57 58 0.5
C9_131 57 193 1.4e-15
C9_132 58 193 1.4e-15
R9_14 44 56 0.35
C9_141 44 193 1.68e-15
C9_142 56 193 1.68e-15
R9_15 43 45 0.2
C9_151 43 193 1.08e-15
C9_152 45 193 1.08e-15
R9_16 46 47 0.5
C9_161 46 193 2.52e-15
C9_162 47 193 2.52e-15
R9_17 45 46 0.05
C9_171 45 193 2.4e-16
C9_172 46 193 2.4e-16
R9_18 53 51 0.15
C9_181 53 193 7.2e-16
C9_182 51 193 7.2e-16
R9_19 47 53 0.05
C9_191 47 193 2.4e-16
C9_192 53 193 2.4e-16
R9_20 50 52 0.15
C9_201 50 193 7.2e-16
C9_202 52 193 7.2e-16
R9_21 41 48 0.2
C9_211 41 193 7e-16
C9_212 48 193 7e-16
R9_22 42 41 0.2
C9_221 42 193 7e-16
C9_222 41 193 7e-16
R9_23 39 42 1
C9_231 39 193 2.8e-15
C9_232 42 193 2.8e-15
R8_1 63 64 0.001
R8_2 70 72 0.001
R8_3 73 72 0.001
R8_4 70 71 0.001
R8_5 75 74 0.001
R8_6 68 67 0.001
R8_7 68 69 600
C8_71 68 193 1.875e-15
C8_72 69 193 1.875e-15
R8_8 66 68 500
C8_81 66 193 1.5e-15
C8_82 68 193 1.5e-15
R8_9 74 77 0.2
C8_91 74 193 7.7e-16
C8_92 77 193 7.7e-16
R8_10 67 74 0.7
C8_101 67 193 2.1e-15
C8_102 74 193 2.1e-15
R8_11 65 67 0.5
C8_111 65 193 1.47e-15
C8_112 67 193 1.47e-15
R8_12 73 75 0.25
C8_121 73 193 1.2e-15
C8_122 75 193 1.2e-15
R8_13 72 76 0.2
C8_131 72 193 7.7e-16
C8_132 76 193 7.7e-16
R8_14 71 72 0.2
C8_141 71 193 7e-16
C8_142 72 193 7e-16
R8_15 64 71 1
C8_151 64 193 2.8e-15
C8_152 71 193 2.8e-15
R7_1 82 81 0.001
R7_2 86 85 0.001
R7_3 86 87 0.001
R7_4 90 89 0.001
R7_5 94 93 0.001
R7_6 98 97 0.001
R7_7 88 98 850
C7_71 88 193 2.625e-15
C7_72 98 193 2.625e-15
R7_8 96 98 150
C7_81 96 193 5.25e-16
C7_82 98 193 5.25e-16
R7_9 97 99 0.2
C7_91 97 193 7.7e-16
C7_92 99 193 7.7e-16
R7_10 93 97 0.5
C7_101 93 193 1.4e-15
C7_102 97 193 1.4e-15
R7_11 95 93 0.5
C7_111 95 193 1.47e-15
C7_112 93 193 1.47e-15
R7_12 89 94 0.6
C7_121 89 193 3e-15
C7_122 94 193 3e-15
R7_13 91 90 0.2
C7_131 91 193 1.08e-15
C7_132 90 193 1.08e-15
R7_14 92 91 0.05
C7_141 92 193 2.4e-16
C7_142 91 193 2.4e-16
R7_15 87 92 0.45
C7_151 87 193 2.28e-15
C7_152 92 193 2.28e-15
R7_16 81 85 1
C7_161 81 193 2.8e-15
C7_162 85 193 2.8e-15
R7_17 83 81 0.5
C7_171 83 193 1.47e-15
C7_172 81 193 1.47e-15
R7_18 82 84 600
C7_181 82 193 1.875e-15
C7_182 84 193 1.875e-15
R7_19 80 82 500
C7_191 80 193 1.5e-15
C7_192 82 193 1.5e-15
R6_1 105 104 0.001
R6_2 108 107 0.001
R6_3 107 109 0.001
R6_4 111 110 0.001
R6_5 113 112 0.001
R6_6 118 117 0.001
R6_7 117 115 0.001
R6_8 116 119 0.001
R6_9 116 122 0.001
R6_10 123 124 0.001
R6_11 122 124 1
C6_111 122 193 2.8e-15
C6_112 124 193 2.8e-15
R6_12 119 122 0.2
C6_121 119 193 7e-16
C6_122 122 193 7e-16
R6_13 115 119 0.2
C6_131 115 193 7e-16
C6_132 119 193 7e-16
R6_14 120 118 0.05
C6_141 120 193 2.4e-16
C6_142 118 193 2.4e-16
R6_15 121 120 0.05
C6_151 121 193 2.4e-16
C6_152 120 193 2.4e-16
R6_16 114 121 0.001
C6_161 114 193 1.2e-16
C6_162 121 193 1.2e-16
R6_17 113 114 0.05
C6_171 113 193 3.6e-16
C6_172 114 193 3.6e-16
R6_18 110 112 0.75
C6_181 110 193 3.6e-15
C6_182 112 193 3.6e-15
R6_19 109 111 0.3
C6_191 109 193 1.44e-15
C6_192 111 193 1.44e-15
R6_20 104 108 1
C6_201 104 193 2.8e-15
C6_202 108 193 2.8e-15
R6_21 103 104 0.2
C6_211 103 193 7.7e-16
C6_212 104 193 7.7e-16
R6_22 105 106 850
C6_221 105 193 2.625e-15
C6_222 106 193 2.625e-15
R6_23 102 105 150
C6_231 102 193 5.25e-16
C6_232 105 193 5.25e-16
R5_1 127 132 0.001
R5_2 129 138 0.001
R5_3 128 137 0.001
R5_4 149 138 0.001
R5_5 148 137 0.001
R5_6 130 139 0.001
R5_7 150 139 0.001
R5_8 131 143 0.001
R5_9 151 143 0.001
R5_10 146 147 0.001
C5_101 146 193 2.145e-15
C5_102 147 193 2.145e-15
R5_11 143 146 0.001
C5_111 143 193 2.34e-15
C5_112 146 193 2.34e-15
R5_12 144 143 0.001
C5_121 144 193 1.365e-15
C5_122 143 193 1.365e-15
R5_13 145 144 0.001
C5_131 145 193 3.9e-16
C5_132 144 193 3.9e-16
R5_14 142 145 0.001
C5_141 142 193 1.755e-15
C5_142 145 193 1.755e-15
R5_15 139 142 0.001
C5_151 139 193 2.34e-15
C5_152 142 193 2.34e-15
R5_16 140 139 0.001
C5_161 140 193 1.365e-15
C5_162 139 193 1.365e-15
R5_17 141 140 0.001
C5_171 141 193 3.9e-16
C5_172 140 193 3.9e-16
R5_18 138 141 0.001
C5_181 138 193 1.365e-15
C5_182 141 193 1.365e-15
R5_19 137 138 0.1
C5_191 137 193 4.7775e-15
C5_192 138 193 4.7775e-15
R5_20 135 137 0.001
C5_201 135 193 1.2675e-15
C5_202 137 193 1.2675e-15
R5_21 136 135 0.001
C5_211 136 193 3.9e-16
C5_212 135 193 3.9e-16
R5_22 134 136 0.001
C5_221 134 193 1.08e-15
C5_222 136 193 1.08e-15
R5_23 132 134 0.1
C5_231 132 193 1.44e-15
C5_232 134 193 1.44e-15
R5_24 133 132 0.001
C5_241 133 193 1.08e-15
C5_242 132 193 1.08e-15
R4_1 154 156 0.001
R4_2 162 163 0.001
R4_3 162 167 0.001
R4_4 164 163 0.001
R4_5 166 165 0.001
R4_6 159 160 0.001
R4_7 159 161 600
C4_71 159 193 1.875e-15
C4_72 161 193 1.875e-15
R4_8 157 159 500
C4_81 157 193 1.5e-15
C4_82 159 193 1.5e-15
R4_9 165 168 0.2
C4_91 165 193 7.7e-16
C4_92 168 193 7.7e-16
R4_10 160 165 0.7
C4_101 160 193 2.1e-15
C4_102 165 193 2.1e-15
R4_11 158 160 0.5
C4_111 158 193 1.47e-15
C4_112 160 193 1.47e-15
R4_12 164 166 0.35
C4_121 164 193 1.8e-15
C4_122 166 193 1.8e-15
R4_13 163 167 0.2
C4_131 163 193 7e-16
C4_132 167 193 7e-16
R4_14 155 163 1.2
C4_141 155 193 3.5e-15
C4_142 163 193 3.5e-15
R4_15 155 156 0.2
C4_151 155 193 5.6e-16
C4_152 156 193 5.6e-16
R3_1 171 172 0.001
R3_2 175 177 0.001
R3_3 181 180 0.001
R3_4 175 178 0.001
R3_5 183 182 0.001
R3_6 176 179 0.001
R3_7 174 176 1150
C3_71 174 193 3.5625e-15
C3_72 176 193 3.5625e-15
R3_8 179 182 0.5
C3_81 179 193 1.4e-15
C3_82 182 193 1.4e-15
R3_9 173 179 1
C3_91 173 193 2.87e-15
C3_92 179 193 2.87e-15
R3_10 181 183 0.25
C3_101 181 193 1.2e-15
C3_102 183 193 1.2e-15
R3_11 177 180 0.2
C3_111 177 193 7e-16
C3_112 180 193 7e-16
R3_12 178 177 0.2
C3_121 178 193 7e-16
C3_122 177 193 7e-16
R3_13 172 178 1
C3_131 172 193 2.8e-15
C3_132 178 193 2.8e-15
R1_1 206 207 0.001
R1_2 211 214 0.001
R1_3 215 216 0.001
R1_4 192 193 0.001
R1_5 197 200 0.001
R1_6 189 190 0.001
R1_7 201 202 0.001
R1_8 202 205 0.1
C1_81 202 193 2.76e-15
C1_82 205 193 2.76e-15
R1_9 203 202 0.001
C1_91 203 193 8.4e-16
C1_92 202 193 8.4e-16
R1_10 190 194 0.1
C1_101 190 193 2.52e-15
C1_102 194 193 2.52e-15
R1_11 191 190 0.001
C1_111 191 193 1.08e-15
C1_112 190 193 1.08e-15
R1_12 204 203 0.001
C1_121 204 193 2.4e-16
C1_122 203 193 2.4e-16
R1_13 200 204 0.1
C1_131 200 193 2.52e-15
C1_132 204 193 2.52e-15
R1_14 198 200 0.001
C1_141 198 193 8.4e-16
C1_142 200 193 8.4e-16
R1_15 199 198 0.001
C1_151 199 193 2.4e-16
C1_152 198 193 2.4e-16
R1_16 196 199 0.1
C1_161 196 193 1.68e-15
C1_162 199 193 1.68e-15
R1_17 193 196 0.1
C1_171 193 193 1.98e-15
C1_172 196 193 1.98e-15
R1_18 195 193 0.001
C1_181 195 193 9e-16
C1_182 193 193 9e-16
R1_19 194 195 0.001
C1_191 194 193 2.4e-16
C1_192 195 193 2.4e-16
R1_20 216 219 0.1
C1_201 216 193 2.76e-15
C1_202 219 193 2.76e-15
R1_21 217 216 0.001
C1_211 217 193 8.4e-16
C1_212 216 193 8.4e-16
R1_22 218 217 0.001
C1_221 218 193 2.4e-16
C1_222 217 193 2.4e-16
R1_23 214 218 0.1
C1_231 214 193 2.52e-15
C1_232 218 193 2.52e-15
R1_24 212 214 0.001
C1_241 212 193 8.4e-16
C1_242 214 193 8.4e-16
R1_25 213 212 0.001
C1_251 213 193 2.4e-16
C1_252 212 193 2.4e-16
R1_26 210 213 0.1
C1_261 210 193 1.68e-15
C1_262 213 193 1.68e-15
R1_27 209 210 0.1
C1_271 209 193 1.56e-15
C1_272 210 193 1.56e-15
R1_28 207 209 0.001
C1_281 207 193 4.8e-16
C1_282 209 193 4.8e-16
R1_29 208 207 0.001
C1_291 208 193 1.08e-15
C1_292 207 193 1.08e-15
.ends 2faseclk

