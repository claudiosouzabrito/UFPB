.include mux4inv.spi

*  d0 d1 d2 d3 s0 s1 vdd vdd2 vss y 
x1 10 11 12 13 14 15 20 20 30 40 mux4inv

r1 40 30 100k

v10 10 30 sine(0.9 0.9 0.25g 0 0 0)
v11 11 30 pulse(0v 1.8v 0s 1ps 8ns 1ps 8ns)
v12 12 30 pulse(0v 1.8v 0s 4ns 4ns 1ps 8ns)
v13 13 30 pulse(0v 1.8v 0s 8ns 1ps 1ps 8ns)

V20 20 30 1.8V
V30 30 0 DC 0
v1 14 30 pulse(0v 1.8v 32ns 1ps 1ps 32ns 64ns)
v2 15 30 pulse(0v 1.8v 16ns 1ps 1ps 16ns 32ns)

.model tp pmos level = 54
.model tn nmos level = 54

.tran 1ps 64ns
.end
