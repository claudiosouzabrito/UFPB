* Spice description of inv+fo4
* Spice driver version -1725303288
* Date ( dd/mm/yyyy hh:mm:ss ): 11/07/2019 at 15:16:11

* INTERF a vdd vss y 


.subckt inv+fo4 29 64 141 85 
* NET 1 = fo4.inv4.inversor_1.nq
* NET 9 = fo4.inv3.inversor_1.nq
* NET 17 = fo4.inv2.inversor_1.nq
* NET 29 = a
* NET 64 = vdd
* NET 85 = y
* NET 108 = fo4.inv1.inversor_1.nq
* NET 141 = vss
Mtr_00020 110 89 35 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00019 35 89 110 64 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00018 19 90 36 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00017 36 90 19 64 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00016 11 95 37 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00015 37 95 11 64 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00014 3 96 38 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00013 38 96 3 64 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00012 99 30 34 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00011 34 30 99 64 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00010 119 70 108 141 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00009 119 70 108 141 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00008 125 71 17 141 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00007 125 71 17 141 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00006 129 74 9 141 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00005 129 74 9 141 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00004 134 75 1 141 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00003 134 75 1 141 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00002 116 26 67 141 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00001 116 26 67 141 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
R8_1 1 2 0.001
R8_2 3 5 0.001
R8_3 3 4 0.001
R8_4 5 6 0.2
C8_41 5 141 7.7e-16
C8_42 6 141 7.7e-16
R8_5 4 5 0.2
C8_51 4 141 7e-16
C8_52 5 141 7e-16
R8_6 2 4 1
C8_61 2 141 2.8e-15
C8_62 4 141 2.8e-15
R7_1 9 10 0.001
R7_2 11 13 0.001
R7_3 11 12 0.001
R7_4 13 14 0.2
C7_41 13 141 7.7e-16
C7_42 14 141 7.7e-16
R7_5 12 13 0.2
C7_51 12 141 7e-16
C7_52 13 141 7e-16
R7_6 10 12 1
C7_61 10 141 2.8e-15
C7_62 12 141 2.8e-15
R6_1 17 18 0.001
R6_2 19 21 0.001
R6_3 19 20 0.001
R6_4 21 22 0.2
C6_41 21 141 7.7e-16
C6_42 22 141 7.7e-16
R6_5 20 21 0.2
C6_51 20 141 7e-16
C6_52 21 141 7e-16
R6_6 18 20 1
C6_61 18 141 2.8e-15
C6_62 20 141 2.8e-15
R5_1 28 27 0.001
R5_2 29 31 0.6
C5_21 29 141 1.75e-15
C5_22 31 141 1.75e-15
R5_3 27 29 0.4
C5_31 27 141 1.12e-15
C5_32 29 141 1.12e-15
R5_4 25 27 0.5
C5_41 25 141 1.47e-15
C5_42 27 141 1.47e-15
R5_5 28 30 700
C5_51 28 141 2.1e-15
C5_52 30 141 2.1e-15
R5_6 26 28 450
C5_61 26 141 1.35e-15
C5_62 28 141 1.35e-15
R4_1 35 45 0.001
R4_2 34 39 0.001
R4_3 36 48 0.001
R4_4 37 53 0.001
R4_5 38 58 0.001
R4_6 61 63 0.001
C4_61 61 141 6e-16
C4_62 63 141 6e-16
R4_7 62 61 0.001
C4_71 62 141 7.2e-16
C4_72 61 141 7.2e-16
R4_8 58 62 0.1
C4_81 58 141 1.56e-15
C4_82 62 141 1.56e-15
R4_9 59 58 0.001
C4_91 59 141 7.2e-16
C4_92 58 141 7.2e-16
R4_10 60 59 0.001
C4_101 60 141 2.4e-16
C4_102 59 141 2.4e-16
R4_11 56 60 0.001
C4_111 56 141 3.6e-16
C4_112 60 141 3.6e-16
R4_12 57 56 0.001
C4_121 57 141 7.2e-16
C4_122 56 141 7.2e-16
R4_13 53 57 0.1
C4_131 53 141 1.56e-15
C4_132 57 141 1.56e-15
R4_14 54 53 0.001
C4_141 54 141 7.2e-16
C4_142 53 141 7.2e-16
R4_15 55 54 0.001
C4_151 55 141 2.4e-16
C4_152 54 141 2.4e-16
R4_16 52 55 0.001
C4_161 52 141 3.6e-16
C4_162 55 141 3.6e-16
R4_17 51 52 0.001
C4_171 51 141 7.2e-16
C4_172 52 141 7.2e-16
R4_18 48 51 0.1
C4_181 48 141 1.56e-15
C4_182 51 141 1.56e-15
R4_19 49 48 0.001
C4_191 49 141 7.2e-16
C4_192 48 141 7.2e-16
R4_20 41 43 0.001
C4_201 41 141 3.6e-16
C4_202 43 141 3.6e-16
R4_21 42 41 0.001
C4_211 42 141 7.2e-16
C4_212 41 141 7.2e-16
R4_22 42 64 0.001
C4_221 42 141 4.8e-16
C4_222 64 141 4.8e-16
R4_23 39 64 0.001
C4_231 39 141 1.08e-15
C4_232 64 141 1.08e-15
R4_24 40 39 0.001
C4_241 40 141 9.6e-16
C4_242 39 141 9.6e-16
R4_25 50 49 0.001
C4_251 50 141 2.4e-16
C4_252 49 141 2.4e-16
R4_26 47 50 0.001
C4_261 47 141 3.6e-16
C4_262 50 141 3.6e-16
R4_27 46 47 0.001
C4_271 46 141 7.2e-16
C4_272 47 141 7.2e-16
R4_28 45 46 0.1
C4_281 45 141 1.56e-15
C4_282 46 141 1.56e-15
R4_29 44 45 0.001
C4_291 44 141 7.2e-16
C4_292 45 141 7.2e-16
R4_30 43 44 0.001
C4_301 43 141 2.4e-16
C4_302 44 141 2.4e-16
R3_1 67 68 0.001
R3_2 99 100 0.001
R3_3 99 85 0.001
R3_4 86 85 0.001
R3_5 88 87 0.001
R3_6 98 97 0.001
R3_7 92 91 0.001
R3_8 94 93 0.001
R3_9 78 77 0.001
R3_10 84 83 0.001
R3_11 80 79 0.001
R3_12 82 81 0.001
R3_13 82 95 700
C3_131 82 141 2.1e-15
C3_132 95 141 2.1e-15
R3_14 74 82 450
C3_141 74 141 1.35e-15
C3_142 82 141 1.35e-15
R3_15 80 90 700
C3_151 80 141 2.1e-15
C3_152 90 141 2.1e-15
R3_16 71 80 450
C3_161 71 141 1.35e-15
C3_162 80 141 1.35e-15
R3_17 84 96 700
C3_171 84 141 2.1e-15
C3_172 96 141 2.1e-15
R3_18 75 84 450
C3_181 75 141 1.35e-15
C3_182 84 141 1.35e-15
R3_19 78 89 700
C3_191 78 141 2.1e-15
C3_192 89 141 2.1e-15
R3_20 70 78 450
C3_201 70 141 1.35e-15
C3_202 78 141 1.35e-15
R3_21 93 104 0.6
C3_211 93 141 1.75e-15
C3_212 104 141 1.75e-15
R3_22 81 93 0.4
C3_221 81 141 1.12e-15
C3_222 93 141 1.12e-15
R3_23 73 81 0.5
C3_231 73 141 1.47e-15
C3_232 81 141 1.47e-15
R3_24 91 103 0.6
C3_241 91 141 1.75e-15
C3_242 103 141 1.75e-15
R3_25 79 91 0.4
C3_251 79 141 1.12e-15
C3_252 91 141 1.12e-15
R3_26 72 79 0.5
C3_261 72 141 1.47e-15
C3_262 79 141 1.47e-15
R3_27 97 105 0.6
C3_271 97 141 1.75e-15
C3_272 105 141 1.75e-15
R3_28 83 97 0.4
C3_281 83 141 1.12e-15
C3_282 97 141 1.12e-15
R3_29 76 83 0.5
C3_291 76 141 1.47e-15
C3_292 83 141 1.47e-15
R3_30 87 102 0.6
C3_301 87 141 1.75e-15
C3_302 102 141 1.75e-15
R3_31 77 87 0.4
C3_311 77 141 1.12e-15
C3_312 87 141 1.12e-15
R3_32 69 77 0.5
C3_321 69 141 1.47e-15
C3_322 77 141 1.47e-15
R3_33 94 98 0.35
C3_331 94 141 1.8e-15
C3_332 98 141 1.8e-15
R3_34 92 94 0.35
C3_341 92 141 1.8e-15
C3_342 94 141 1.8e-15
R3_35 88 92 0.35
C3_351 88 141 1.8e-15
C3_352 92 141 1.8e-15
R3_36 86 88 0.25
C3_361 86 141 1.2e-15
C3_362 88 141 1.2e-15
R3_37 100 101 0.2
C3_371 100 141 7.7e-16
C3_372 101 141 7.7e-16
R3_38 85 100 0.3
C3_381 85 141 8.4e-16
C3_382 100 141 8.4e-16
R3_39 68 85 0.9
C3_391 68 141 2.66e-15
C3_392 85 141 2.66e-15
R2_1 108 109 0.001
R2_2 110 112 0.001
R2_3 110 111 0.001
R2_4 112 113 0.2
C2_41 112 141 7.7e-16
C2_42 113 141 7.7e-16
R2_5 111 112 0.2
C2_51 111 141 7e-16
C2_52 112 141 7e-16
R2_6 109 111 1
C2_61 109 141 2.8e-15
C2_62 111 141 2.8e-15
R1_1 119 120 0.001
R1_2 116 117 0.001
R1_3 125 126 0.001
R1_4 129 131 0.001
R1_5 134 136 0.001
R1_6 139 140 0.001
C1_61 139 141 6e-16
C1_62 140 141 6e-16
R1_7 136 139 0.1
C1_71 136 141 2.28e-15
C1_72 139 141 2.28e-15
R1_8 137 136 0.001
C1_81 137 141 7.2e-16
C1_82 136 141 7.2e-16
R1_9 138 137 0.001
C1_91 138 141 2.4e-16
C1_92 137 141 2.4e-16
R1_10 135 138 0.001
C1_101 135 141 3.6e-16
C1_102 138 141 3.6e-16
R1_11 131 135 0.1
C1_111 131 141 2.28e-15
C1_112 135 141 2.28e-15
R1_12 132 131 0.001
C1_121 132 141 7.2e-16
C1_122 131 141 7.2e-16
R1_13 133 132 0.001
C1_131 133 141 2.4e-16
C1_132 132 141 2.4e-16
R1_14 130 133 0.001
C1_141 130 141 3.6e-16
C1_142 133 141 3.6e-16
R1_15 126 130 0.1
C1_151 126 141 2.28e-15
C1_152 130 141 2.28e-15
R1_16 127 126 0.001
C1_161 127 141 7.2e-16
C1_162 126 141 7.2e-16
R1_17 121 122 0.001
C1_171 121 141 3.6e-16
C1_172 122 141 3.6e-16
R1_18 121 141 0.001
C1_181 121 141 1.2e-15
C1_182 141 141 1.2e-15
R1_19 117 141 0.001
C1_191 117 141 1.08e-15
C1_192 141 141 1.08e-15
R1_20 118 117 0.001
C1_201 118 141 9.6e-16
C1_202 117 141 9.6e-16
R1_21 128 127 0.001
C1_211 128 141 2.4e-16
C1_212 127 141 2.4e-16
R1_22 124 128 0.001
C1_221 124 141 3.6e-16
C1_222 128 141 3.6e-16
R1_23 120 124 0.1
C1_231 120 141 2.28e-15
C1_232 124 141 2.28e-15
R1_24 123 120 0.001
C1_241 123 141 7.2e-16
C1_242 120 141 7.2e-16
R1_25 122 123 0.001
C1_251 122 141 2.4e-16
C1_252 123 141 2.4e-16
.ends inv+fo4

