.include biel10.spi

x1 10 20 30 40 42 44 biel10

V1 20 30 1.8V
V2 10 30 0V DC
V3 30 0 DC 0

.model tp pmos level = 54
.model tn nmos level = 54

.dc V2 0 1.8 0.001
.end
