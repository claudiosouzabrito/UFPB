* Spice description of inversor4
* Spice driver version 341243400
* Date ( dd/mm/yyyy hh:mm:ss ): 30/06/2019 at 15:24:36

* INTERF a vdd vss y 


.subckt inversor4 5 16 31 22 
* NET 5 = a
* NET 16 = vdd
* NET 22 = y
* NET 31 = vss
Mtr_00004 21 6 10 16 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00003 10 6 21 16 tp L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00002 28 2 19 31 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00001 28 2 19 31 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
R4_1 4 3 0.001
R4_2 5 7 0.6
C4_21 5 31 1.75e-15
C4_22 7 31 1.75e-15
R4_3 3 5 0.4
C4_31 3 31 1.12e-15
C4_32 5 31 1.12e-15
R4_4 1 3 0.5
C4_41 1 31 1.47e-15
C4_42 3 31 1.47e-15
R4_5 4 6 700
C4_51 4 31 2.1e-15
C4_52 6 31 2.1e-15
R4_6 2 4 450
C4_61 2 31 1.35e-15
C4_62 4 31 1.35e-15
R3_1 10 11 0.001
R3_2 14 15 0.001
C3_21 14 31 6e-16
C3_22 15 31 6e-16
R3_3 13 14 0.001
C3_31 13 31 7.2e-16
C3_32 14 31 7.2e-16
R3_4 13 16 0.001
C3_41 13 31 4.8e-16
C3_42 16 31 4.8e-16
R3_5 11 16 0.001
C3_51 11 31 1.08e-15
C3_52 16 31 1.08e-15
R3_6 12 11 0.001
C3_61 12 31 9.6e-16
C3_62 11 31 9.6e-16
R2_1 19 20 0.001
R2_2 21 24 0.001
R2_3 21 23 0.001
R2_4 24 25 0.2
C2_41 24 31 7.7e-16
C2_42 25 31 7.7e-16
R2_5 23 24 0.2
C2_51 23 31 7e-16
C2_52 24 31 7e-16
R2_6 22 23 0.1
C2_61 22 31 2.8e-16
C2_62 23 31 2.8e-16
R2_7 20 22 0.9
C2_71 20 31 2.52e-15
C2_72 22 31 2.52e-15
R1_1 28 29 0.001
R1_2 32 33 0.001
C1_21 32 31 6e-16
C1_22 33 31 6e-16
R1_3 32 31 0.001
C1_31 32 31 1.2e-15
C1_32 31 31 1.2e-15
R1_4 29 31 0.001
C1_41 29 31 1.08e-15
C1_42 31 31 1.08e-15
R1_5 30 29 0.001
C1_51 30 31 9.6e-16
C1_52 29 31 9.6e-16
.ends inversor4

