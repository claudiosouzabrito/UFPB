* Spice description of nand2
* Spice driver version 1093072392
* Date ( dd/mm/yyyy hh:mm:ss ): 25/07/2019 at 15:22:51

* INTERF a0 a1 vdd vss y 


.subckt nand2 5 47 19 23 36 
* NET 5 = a0
* NET 19 = vdd
* NET 23 = vss
* NET 36 = y
* NET 47 = a1
Mtr_00006 34 6 10 19 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00005 34 48 11 19 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00004 10 6 34 19 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00003 22 2 32 23 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00002 32 42 41 23 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00001 22 2 32 23 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
R5_1 4 3 0.001
R5_2 5 7 0.6
C5_21 5 23 1.89e-15
C5_22 7 23 1.89e-15
R5_3 3 5 0.3
C5_31 3 23 9.8e-16
C5_32 5 23 9.8e-16
R5_4 1 3 0.5
C5_41 1 23 1.47e-15
C5_42 3 23 1.47e-15
R5_5 4 6 700
C5_51 4 23 2.1e-15
C5_52 6 23 2.1e-15
R5_6 2 4 450
C5_61 2 23 1.35e-15
C5_62 4 23 1.35e-15
R4_1 10 12 0.001
R4_2 10 13 0.001
R4_3 11 17 0.001
R4_4 17 18 0.001
C4_41 17 23 8.4e-16
C4_42 18 23 8.4e-16
R4_5 16 17 0.1
C4_51 16 23 1.56e-15
C4_52 17 23 1.56e-15
R4_6 15 16 0.001
C4_61 15 23 1.2e-15
C4_62 16 23 1.2e-15
R4_7 15 19 0.001
C4_71 15 23 1.08e-15
C4_72 19 23 1.08e-15
R4_8 13 19 0.001
C4_81 13 23 4.8e-16
C4_82 19 23 4.8e-16
R4_9 12 13 0.001
C4_91 12 23 7.2e-16
C4_92 13 23 7.2e-16
R4_10 14 12 0.001
C4_101 14 23 3.6e-16
C4_102 12 23 3.6e-16
R3_1 22 24 0.001
R3_2 22 25 0.001
R3_3 28 29 0.1
C3_31 28 23 2.4e-15
C3_32 29 23 2.4e-15
R3_4 27 28 0.001
C3_41 27 23 1.08e-15
C3_42 28 23 1.08e-15
R3_5 27 23 0.001
C3_51 27 23 1.2e-15
C3_52 23 23 1.2e-15
R3_6 25 23 0.001
C3_61 25 23 4.8e-16
C3_62 23 23 4.8e-16
R3_7 24 25 0.001
C3_71 24 23 7.2e-16
C3_72 25 23 7.2e-16
R3_8 26 24 0.001
C3_81 26 23 3.6e-16
C3_82 24 23 3.6e-16
R2_1 32 33 0.001
R2_2 34 37 0.001
R2_3 34 35 0.001
R2_4 37 38 0.2
C2_41 37 23 7.7e-16
C2_42 38 23 7.7e-16
R2_5 35 37 0.2
C2_51 35 23 7e-16
C2_52 37 23 7e-16
R2_6 36 35 0.1
C2_61 36 23 2.8e-16
C2_62 35 23 2.8e-16
R2_7 33 36 0.9
C2_71 33 23 2.52e-15
C2_72 36 23 2.52e-15
R1_1 41 43 0.001
R1_2 50 49 0.001
R1_3 50 48 650
C1_31 50 23 1.95e-15
C1_32 48 23 1.95e-15
R1_4 42 50 450
C1_41 42 23 1.35e-15
C1_42 50 23 1.35e-15
R1_5 47 51 0.6
C1_51 47 23 1.89e-15
C1_52 51 23 1.89e-15
R1_6 49 47 0.3
C1_61 49 23 8.4e-16
C1_62 47 23 8.4e-16
R1_7 44 49 0.2
C1_71 44 23 6.3e-16
C1_72 49 23 6.3e-16
R1_8 45 44 0.001
C1_81 45 23 1.4e-16
C1_82 44 23 1.4e-16
R1_9 43 45 0.2
C1_91 43 23 6.3e-16
C1_92 45 23 6.3e-16
R1_10 46 43 0.001
C1_101 46 23 2.1e-16
C1_102 43 23 2.1e-16
.ends nand2

