* Spice description of mux4inv
* Spice driver version -1024231928
* Date ( dd/mm/yyyy hh:mm:ss ):  6/08/2019 at 15:31:30

* INTERF d0 d1 d2 d3 s0 s1 vdd vdd2 vss y 


.subckt mux4inv 214 182 389 360 477 150 59 503 329 76 
* NET 59 = vdd
* NET 76 = y
* NET 91 = mux3.tirs2.inversor_1.nq
* NET 109 = mux3.tirs1.inversor_1.nq
* NET 150 = s1
* NET 157 = mux3.inv1.inversor_1.nq
* NET 182 = d1
* NET 193 = mux1.tirs2.inversor_1.nq
* NET 214 = d0
* NET 263 = mux1.inv1.inversor_1.nq
* NET 288 = mux1.tirs1.inversor_1.nq
* NET 329 = vss
* NET 360 = d3
* NET 369 = mux2.tirs2.inversor_1.nq
* NET 389 = d2
* NET 477 = s0
* NET 485 = mux2.tirs1.inversor_1.nq
* NET 503 = vdd2
* NET 529 = mux2.inv1.inversor_1.nq
Mtr_00066 96 152 21 503 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00065 22 423 1 503 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00064 1 98 77 503 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00063 21 152 96 503 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00062 114 176 19 503 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00061 20 239 4 503 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00060 4 116 73 503 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00059 19 176 114 503 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00058 172 149 18 503 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00057 18 149 172 503 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00056 369 435 517 503 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00055 524 359 366 503 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00054 366 374 401 503 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00053 517 435 369 503 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00052 485 532 509 503 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00051 514 388 430 503 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00050 430 490 395 503 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00049 509 532 485 503 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00048 529 433 504 503 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00047 504 433 529 503 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00046 198 480 16 503 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00045 17 187 7 503 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00044 7 200 242 503 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00043 16 480 198 503 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00042 293 282 13 503 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00041 15 219 10 503 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00040 10 295 240 503 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00039 13 282 293 503 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00038 278 478 14 503 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00037 14 478 278 503 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00036 355 132 91 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00035 346 420 62 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00034 62 138 69 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00033 355 132 91 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00032 62 138 69 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00031 354 160 109 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00030 339 230 127 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00029 127 165 65 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00028 354 160 109 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00027 127 165 65 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00026 353 130 157 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00025 353 130 157 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00024 309 447 383 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00023 310 363 211 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00022 211 450 415 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00021 309 447 383 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00020 211 450 415 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00019 306 540 499 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00018 308 392 260 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00017 260 541 411 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00016 306 540 499 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00015 260 541 411 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00014 307 444 542 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00013 307 444 542 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00012 352 459 193 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00011 331 185 190 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00010 190 471 226 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00009 352 459 193 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00008 190 471 226 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00007 350 266 288 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00006 330 217 257 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00005 257 271 222 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00004 350 266 288 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00003 257 271 222 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00002 351 458 263 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00001 351 458 263 329 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
R29_1 13 23 0.001
R29_2 15 32 0.001
R29_3 17 39 0.001
R29_4 16 33 0.001
R29_5 14 25 0.001
R29_6 18 40 0.001
R29_7 20 49 0.001
R29_8 19 46 0.001
R29_9 22 55 0.001
R29_10 21 51 0.001
R29_11 55 58 0.3
C29_111 55 329 4.92e-15
C29_112 58 329 4.92e-15
R29_12 57 55 0.1
C29_121 57 329 2.28e-15
C29_122 55 329 2.28e-15
R29_13 56 57 0.001
C29_131 56 329 1.32e-15
C29_132 57 329 1.32e-15
R29_14 51 56 0.1
C29_141 51 329 1.56e-15
C29_142 56 329 1.56e-15
R29_15 52 51 0.001
C29_151 52 329 7.2e-16
C29_152 51 329 7.2e-16
R29_16 53 52 0.001
C29_161 53 329 2.4e-16
C29_162 52 329 2.4e-16
R29_17 54 53 0.001
C29_171 54 329 2.4e-16
C29_172 53 329 2.4e-16
R29_18 49 54 0.3
C29_181 49 329 4.44e-15
C29_182 54 329 4.44e-15
R29_19 50 49 0.1
C29_191 50 329 2.28e-15
C29_192 49 329 2.28e-15
R29_20 45 50 0.001
C29_201 45 329 1.32e-15
C29_202 50 329 1.32e-15
R29_21 46 45 0.1
C29_211 46 329 1.56e-15
C29_212 45 329 1.56e-15
R29_22 47 46 0.001
C29_221 47 329 7.2e-16
C29_222 46 329 7.2e-16
R29_23 48 47 0.001
C29_231 48 329 2.4e-16
C29_232 47 329 2.4e-16
R29_24 43 48 0.001
C29_241 43 329 3.6e-16
C29_242 48 329 3.6e-16
R29_25 44 43 0.001
C29_251 44 329 7.2e-16
C29_252 43 329 7.2e-16
R29_26 40 44 0.1
C29_261 40 329 1.56e-15
C29_262 44 329 1.56e-15
R29_27 41 40 0.001
C29_271 41 329 7.2e-16
C29_272 40 329 7.2e-16
R29_28 26 24 0.001
C29_281 26 329 7.2e-16
C29_282 24 329 7.2e-16
R29_29 26 59 0.001
C29_291 26 329 4.8e-16
C29_292 59 329 4.8e-16
R29_30 25 59 0.001
C29_301 25 329 1.08e-15
C29_302 59 329 1.08e-15
R29_31 29 25 0.001
C29_311 29 329 9.6e-16
C29_312 25 329 9.6e-16
R29_32 42 41 0.001
C29_321 42 329 2.4e-16
C29_322 41 329 2.4e-16
R29_33 39 42 0.3
C29_331 39 329 4.68e-15
C29_332 42 329 4.68e-15
R29_34 36 39 0.1
C29_341 36 329 2.28e-15
C29_342 39 329 2.28e-15
R29_35 34 36 0.001
C29_351 34 329 1.32e-15
C29_352 36 329 1.32e-15
R29_36 33 34 0.1
C29_361 33 329 1.56e-15
C29_362 34 329 1.56e-15
R29_37 35 33 0.001
C29_371 35 329 7.2e-16
C29_372 33 329 7.2e-16
R29_38 37 35 0.001
C29_381 37 329 2.4e-16
C29_382 35 329 2.4e-16
R29_39 38 37 0.001
C29_391 38 329 2.4e-16
C29_392 37 329 2.4e-16
R29_40 32 38 0.3
C29_401 32 329 4.44e-15
C29_402 38 329 4.44e-15
R29_41 31 32 0.1
C29_411 31 329 2.28e-15
C29_412 32 329 2.28e-15
R29_42 30 31 0.001
C29_421 30 329 1.32e-15
C29_422 31 329 1.32e-15
R29_43 23 30 0.1
C29_431 23 329 1.56e-15
C29_432 30 329 1.56e-15
R29_44 28 23 0.001
C29_441 28 329 7.2e-16
C29_442 23 329 7.2e-16
R29_45 27 28 0.001
C29_451 27 329 2.4e-16
C29_452 28 329 2.4e-16
R29_46 24 27 0.001
C29_461 24 329 3.6e-16
C29_462 27 329 3.6e-16
R27_1 65 66 0.001
R27_2 75 74 0.001
R27_3 73 83 0.001
R27_4 78 76 0.001
R27_5 77 86 0.001
R27_6 69 70 0.001
R27_7 70 71 0.1
C27_71 70 329 1.725e-16
C27_72 71 329 1.725e-16
R27_8 86 88 0.2
C27_81 86 329 2.875e-16
C27_82 88 329 2.875e-16
R27_9 87 86 0.1
C27_91 87 329 1.725e-16
C27_92 86 329 1.725e-16
R27_10 81 87 0.1
C27_101 81 329 1.15e-16
C27_102 87 329 1.15e-16
R27_11 76 81 1
C27_111 76 329 1.2075e-15
C27_112 81 329 1.2075e-15
R27_12 72 76 0.9
C27_121 72 329 1.0925e-15
C27_122 76 329 1.0925e-15
R27_13 71 72 0.1
C27_131 71 329 1.15e-16
C27_132 72 329 1.15e-16
R27_14 78 82 0.15
C27_141 78 329 8.4e-16
C27_142 82 329 8.4e-16
R27_15 79 82 1.1
C27_151 79 329 5.4e-15
C27_152 82 329 5.4e-15
R27_16 75 79 0.15
C27_161 75 329 8.4e-16
C27_162 79 329 8.4e-16
R27_17 83 85 0.2
C27_171 83 329 2.875e-16
C27_172 85 329 2.875e-16
R27_18 84 83 0.1
C27_181 84 329 1.725e-16
C27_182 83 329 1.725e-16
R27_19 80 84 0.1
C27_191 80 329 1.15e-16
C27_192 84 329 1.15e-16
R27_20 74 80 1
C27_201 74 329 1.2075e-15
C27_202 80 329 1.2075e-15
R27_21 67 74 0.9
C27_211 67 329 1.0925e-15
C27_212 74 329 1.0925e-15
R27_22 68 67 0.1
C27_221 68 329 1.15e-16
C27_222 67 329 1.15e-16
R27_23 66 68 0.1
C27_231 66 329 1.725e-16
C27_232 68 329 1.725e-16
R26_1 91 92 0.001
R26_2 94 93 0.001
R26_3 96 99 0.001
R26_4 96 97 0.001
R26_5 98 104 400
C26_51 98 329 1.275e-15
C26_52 104 329 1.275e-15
R26_6 105 106 50
C26_61 105 329 2.25e-16
C26_62 106 329 2.25e-16
R26_7 104 105 50
C26_71 104 329 1.5e-16
C26_72 105 329 1.5e-16
R26_8 102 106 700
C26_81 102 329 2.175e-15
C26_82 106 329 2.175e-15
R26_9 103 102 50
C26_91 103 329 1.5e-16
C26_92 102 329 1.5e-16
R26_10 101 103 300
C26_101 101 329 9.75e-16
C26_102 103 329 9.75e-16
R26_11 95 101 1200
C26_111 95 329 3.6e-15
C26_112 101 329 3.6e-15
R26_12 94 95 200
C26_121 94 329 6e-16
C26_122 95 329 6e-16
R26_13 99 100 0.2
C26_131 99 329 7.7e-16
C26_132 100 329 7.7e-16
R26_14 97 99 0.2
C26_141 97 329 7e-16
C26_142 99 329 7e-16
R26_15 93 97 0.5
C26_151 93 329 1.4e-15
C26_152 97 329 1.4e-15
R26_16 92 93 0.5
C26_161 92 329 1.4e-15
C26_162 93 329 1.4e-15
R25_1 109 110 0.001
R25_2 112 111 0.001
R25_3 114 117 0.001
R25_4 114 115 0.001
R25_5 116 122 400
C25_51 116 329 1.275e-15
C25_52 122 329 1.275e-15
R25_6 123 124 50
C25_61 123 329 2.25e-16
C25_62 124 329 2.25e-16
R25_7 122 123 50
C25_71 122 329 1.5e-16
C25_72 123 329 1.5e-16
R25_8 120 124 700
C25_81 120 329 2.175e-15
C25_82 124 329 2.175e-15
R25_9 121 120 50
C25_91 121 329 1.5e-16
C25_92 120 329 1.5e-16
R25_10 119 121 300
C25_101 119 329 9.75e-16
C25_102 121 329 9.75e-16
R25_11 113 119 1200
C25_111 113 329 3.6e-15
C25_112 119 329 3.6e-15
R25_12 112 113 200
C25_121 112 329 6e-16
C25_122 113 329 6e-16
R25_13 117 118 0.2
C25_131 117 329 7.7e-16
C25_132 118 329 7.7e-16
R25_14 115 117 0.2
C25_141 115 329 7e-16
C25_142 117 329 7e-16
R25_15 111 115 0.5
C25_151 111 329 1.4e-15
C25_152 115 329 1.4e-15
R25_16 110 111 0.5
C25_161 110 329 1.4e-15
C25_162 111 329 1.4e-15
R23_1 145 144 0.001
R23_2 151 150 0.001
R23_3 147 146 0.001
R23_4 146 148 0.001
R23_5 139 138 200
C23_51 139 329 6.75e-16
C23_52 138 329 6.75e-16
R23_6 140 139 50
C23_61 140 329 1.5e-16
C23_62 139 329 1.5e-16
R23_7 141 140 50
C23_71 141 329 2.25e-16
C23_72 140 329 2.25e-16
R23_8 134 141 700
C23_81 134 329 2.175e-15
C23_82 141 329 2.175e-15
R23_9 135 134 50
C23_91 135 329 1.5e-16
C23_92 134 329 1.5e-16
R23_10 136 135 300
C23_101 136 329 9.75e-16
C23_102 135 329 9.75e-16
R23_11 136 137 100
C23_111 136 329 3e-16
C23_112 137 329 3e-16
R23_12 132 137 400
C23_121 132 329 1.2e-15
C23_122 137 329 1.2e-15
R23_13 148 152 700
C23_131 148 329 2.1e-15
C23_132 152 329 2.1e-15
R23_14 132 148 450
C23_141 132 329 1.35e-15
C23_142 148 329 1.35e-15
R23_15 146 154 1
C23_151 146 329 2.87e-15
C23_152 154 329 2.87e-15
R23_16 133 146 0.5
C23_161 133 329 1.47e-15
C23_162 146 329 1.47e-15
R23_17 143 147 0.1
C23_171 143 329 6e-16
C23_172 147 329 6e-16
R23_18 142 143 1.5
C23_181 142 329 7.2e-15
C23_182 143 329 7.2e-15
R23_19 142 151 0.3
C23_191 142 329 1.56e-15
C23_192 151 329 1.56e-15
R23_20 150 153 0.6
C23_201 150 329 1.75e-15
C23_202 153 329 1.75e-15
R23_21 144 150 0.4
C23_211 144 329 1.12e-15
C23_212 150 329 1.12e-15
R23_22 131 144 0.5
C23_221 131 329 1.47e-15
C23_222 144 329 1.47e-15
R23_23 145 149 700
C23_231 145 329 2.1e-15
C23_232 149 329 2.1e-15
R23_24 130 145 450
C23_241 130 329 1.35e-15
C23_242 145 329 1.35e-15
R22_1 157 158 0.001
R22_2 172 177 0.001
R22_3 172 173 0.001
R22_4 174 173 0.001
R22_5 170 169 0.001
R22_6 169 171 0.001
R22_7 166 165 200
C22_71 166 329 6.75e-16
C22_72 165 329 6.75e-16
R22_8 167 166 50
C22_81 167 329 1.5e-16
C22_82 166 329 1.5e-16
R22_9 168 167 50
C22_91 168 329 2.25e-16
C22_92 167 329 2.25e-16
R22_10 163 168 700
C22_101 163 329 2.175e-15
C22_102 168 329 2.175e-15
R22_11 164 163 50
C22_111 164 329 1.5e-16
C22_112 163 329 1.5e-16
R22_12 161 164 300
C22_121 161 329 9.75e-16
C22_122 164 329 9.75e-16
R22_13 161 162 100
C22_131 161 329 3e-16
C22_132 162 329 3e-16
R22_14 160 162 400
C22_141 160 329 1.2e-15
C22_142 162 329 1.2e-15
R22_15 171 176 700
C22_151 171 329 2.1e-15
C22_152 176 329 2.1e-15
R22_16 160 171 450
C22_161 160 329 1.35e-15
C22_162 171 329 1.35e-15
R22_17 169 179 1
C22_171 169 329 2.87e-15
C22_172 179 329 2.87e-15
R22_18 159 169 0.5
C22_181 159 329 1.47e-15
C22_182 169 329 1.47e-15
R22_19 170 175 0.2
C22_191 170 329 9.6e-16
C22_192 175 329 9.6e-16
R22_20 174 175 0.25
C22_201 174 329 1.2e-15
C22_202 175 329 1.2e-15
R22_21 177 178 0.2
C22_211 177 329 7.7e-16
C22_212 178 329 7.7e-16
R22_22 173 177 0.3
C22_221 173 329 8.4e-16
C22_222 177 329 8.4e-16
R22_23 158 173 0.9
C22_231 158 329 2.66e-15
C22_232 173 329 2.66e-15
R21_1 183 182 0.001
R21_2 182 186 1.5
C21_21 182 329 1.7825e-15
C21_22 186 329 1.7825e-15
R21_3 184 182 0.9
C21_31 184 329 1.0925e-15
C21_32 182 329 1.0925e-15
R21_4 183 187 550
C21_41 183 329 1.65e-15
C21_42 187 329 1.65e-15
R21_5 185 183 500
C21_51 185 329 1.5e-15
C21_52 183 329 1.5e-15
R19_1 193 194 0.001
R19_2 196 195 0.001
R19_3 198 201 0.001
R19_4 198 199 0.001
R19_5 200 206 400
C19_51 200 329 1.275e-15
C19_52 206 329 1.275e-15
R19_6 207 208 50
C19_61 207 329 2.25e-16
C19_62 208 329 2.25e-16
R19_7 206 207 50
C19_71 206 329 1.5e-16
C19_72 207 329 1.5e-16
R19_8 204 208 700
C19_81 204 329 2.175e-15
C19_82 208 329 2.175e-15
R19_9 205 204 50
C19_91 205 329 1.5e-16
C19_92 204 329 1.5e-16
R19_10 203 205 300
C19_101 203 329 9.75e-16
C19_102 205 329 9.75e-16
R19_11 197 203 1200
C19_111 197 329 3.6e-15
C19_112 203 329 3.6e-15
R19_12 196 197 200
C19_121 196 329 6e-16
C19_122 197 329 6e-16
R19_13 201 202 0.2
C19_131 201 329 7.7e-16
C19_132 202 329 7.7e-16
R19_14 199 201 0.2
C19_141 199 329 7e-16
C19_142 201 329 7e-16
R19_15 195 199 0.5
C19_151 195 329 1.4e-15
C19_152 199 329 1.4e-15
R19_16 194 195 0.5
C19_161 194 329 1.4e-15
C19_162 195 329 1.4e-15
R17_1 215 214 0.001
R17_2 214 218 1.5
C17_21 214 329 1.7825e-15
C17_22 218 329 1.7825e-15
R17_3 216 214 0.9
C17_31 216 329 1.0925e-15
C17_32 214 329 1.0925e-15
R17_4 215 219 550
C17_41 215 329 1.65e-15
C17_42 219 329 1.65e-15
R17_5 217 215 500
C17_51 217 329 1.5e-15
C17_52 215 329 1.5e-15
R16_1 222 223 0.001
R16_2 233 232 0.001
R16_3 240 244 0.001
R16_4 235 234 0.001
R16_5 237 236 0.001
R16_6 226 227 0.001
R16_7 242 247 0.001
R16_8 236 238 0.001
R16_9 238 239 550
C16_91 238 329 1.65e-15
C16_92 239 329 1.65e-15
R16_10 230 238 500
C16_101 230 329 1.5e-15
C16_102 238 329 1.5e-15
R16_11 236 254 1.5
C16_111 236 329 1.7825e-15
C16_112 254 329 1.7825e-15
R16_12 231 236 0.9
C16_121 231 329 1.0925e-15
C16_122 236 329 1.0925e-15
R16_13 247 253 0.2
C16_131 247 329 2.875e-16
C16_132 253 329 2.875e-16
R16_14 248 247 0.1
C16_141 248 329 1.725e-16
C16_142 247 329 1.725e-16
R16_15 227 228 0.1
C16_151 227 329 1.725e-16
C16_152 228 329 1.725e-16
R16_16 237 251 0.35
C16_161 237 329 1.68e-15
C16_162 251 329 1.68e-15
R16_17 249 248 0.1
C16_171 249 329 1.15e-16
C16_172 248 329 1.15e-16
R16_18 234 249 1
C16_181 234 329 1.2075e-15
C16_182 249 329 1.2075e-15
R16_19 229 234 0.9
C16_191 229 329 1.0925e-15
C16_192 234 329 1.0925e-15
R16_20 228 229 0.1
C16_201 228 329 1.15e-16
C16_202 229 329 1.15e-16
R16_21 250 251 1.15
C16_211 250 329 5.64e-15
C16_212 251 329 5.64e-15
R16_22 243 250 0.15
C16_221 243 329 8.4e-16
C16_222 250 329 8.4e-16
R16_23 235 243 0.15
C16_231 235 329 8.4e-16
C16_232 243 329 8.4e-16
R16_24 241 243 1.1
C16_241 241 329 5.4e-15
C16_242 243 329 5.4e-15
R16_25 233 241 0.15
C16_251 233 329 8.4e-16
C16_252 241 329 8.4e-16
R16_26 244 252 0.2
C16_261 244 329 2.875e-16
C16_262 252 329 2.875e-16
R16_27 245 244 0.1
C16_271 245 329 1.725e-16
C16_272 244 329 1.725e-16
R16_28 246 245 0.1
C16_281 246 329 1.15e-16
C16_282 245 329 1.15e-16
R16_29 232 246 1
C16_291 232 329 1.2075e-15
C16_292 246 329 1.2075e-15
R16_30 224 232 0.9
C16_301 224 329 1.0925e-15
C16_302 232 329 1.0925e-15
R16_31 225 224 0.1
C16_311 225 329 1.15e-16
C16_312 224 329 1.15e-16
R16_32 223 225 0.1
C16_321 223 329 1.725e-16
C16_322 225 329 1.725e-16
R13_1 263 264 0.001
R13_2 278 283 0.001
R13_3 278 279 0.001
R13_4 280 279 0.001
R13_5 276 275 0.001
R13_6 275 277 0.001
R13_7 272 271 200
C13_71 272 329 6.75e-16
C13_72 271 329 6.75e-16
R13_8 273 272 50
C13_81 273 329 1.5e-16
C13_82 272 329 1.5e-16
R13_9 274 273 50
C13_91 274 329 2.25e-16
C13_92 273 329 2.25e-16
R13_10 269 274 700
C13_101 269 329 2.175e-15
C13_102 274 329 2.175e-15
R13_11 270 269 50
C13_111 270 329 1.5e-16
C13_112 269 329 1.5e-16
R13_12 267 270 300
C13_121 267 329 9.75e-16
C13_122 270 329 9.75e-16
R13_13 267 268 100
C13_131 267 329 3e-16
C13_132 268 329 3e-16
R13_14 266 268 400
C13_141 266 329 1.2e-15
C13_142 268 329 1.2e-15
R13_15 277 282 700
C13_151 277 329 2.1e-15
C13_152 282 329 2.1e-15
R13_16 266 277 450
C13_161 266 329 1.35e-15
C13_162 277 329 1.35e-15
R13_17 275 285 1
C13_171 275 329 2.87e-15
C13_172 285 329 2.87e-15
R13_18 265 275 0.5
C13_181 265 329 1.47e-15
C13_182 275 329 1.47e-15
R13_19 276 281 0.2
C13_191 276 329 9.6e-16
C13_192 281 329 9.6e-16
R13_20 280 281 0.25
C13_201 280 329 1.2e-15
C13_202 281 329 1.2e-15
R13_21 283 284 0.2
C13_211 283 329 7.7e-16
C13_212 284 329 7.7e-16
R13_22 279 283 0.3
C13_221 279 329 8.4e-16
C13_222 283 329 8.4e-16
R13_23 264 279 0.9
C13_231 264 329 2.66e-15
C13_232 279 329 2.66e-15
R12_1 288 289 0.001
R12_2 293 294 0.001
R12_3 293 296 0.001
R12_4 291 290 0.001
R12_5 295 301 400
C12_51 295 329 1.275e-15
C12_52 301 329 1.275e-15
R12_6 302 303 50
C12_61 302 329 2.25e-16
C12_62 303 329 2.25e-16
R12_7 301 302 50
C12_71 301 329 1.5e-16
C12_72 302 329 1.5e-16
R12_8 299 303 700
C12_81 299 329 2.175e-15
C12_82 303 329 2.175e-15
R12_9 300 299 50
C12_91 300 329 1.5e-16
C12_92 299 329 1.5e-16
R12_10 298 300 300
C12_101 298 329 9.75e-16
C12_102 300 329 9.75e-16
R12_11 292 298 1200
C12_111 292 329 3.6e-15
C12_112 298 329 3.6e-15
R12_12 291 292 200
C12_121 291 329 6e-16
C12_122 292 329 6e-16
R12_13 296 297 0.2
C12_131 296 329 7.7e-16
C12_132 297 329 7.7e-16
R12_14 294 296 0.2
C12_141 294 329 7e-16
C12_142 296 329 7e-16
R12_15 290 294 0.5
C12_151 290 329 1.4e-15
C12_152 294 329 1.4e-15
R12_16 289 290 0.5
C12_161 289 329 1.4e-15
C12_162 290 329 1.4e-15
R11_1 306 311 0.001
R11_2 308 319 0.001
R11_3 307 313 0.001
R11_4 330 319 0.001
R11_5 350 311 0.001
R11_6 351 313 0.001
R11_7 309 321 0.001
R11_8 331 325 0.001
R11_9 352 321 0.001
R11_10 310 325 0.001
R11_11 353 333 0.001
R11_12 339 340 0.001
R11_13 354 334 0.001
R11_14 346 347 0.001
R11_15 355 341 0.001
R11_16 347 349 0.3
C11_161 347 329 4.92e-15
C11_162 349 329 4.92e-15
R11_17 348 347 0.1
C11_171 348 329 2.28e-15
C11_172 347 329 2.28e-15
R11_18 342 348 0.001
C11_181 342 329 1.32e-15
C11_182 348 329 1.32e-15
R11_19 341 342 0.1
C11_191 341 329 1.56e-15
C11_192 342 329 1.56e-15
R11_20 343 341 0.001
C11_201 343 329 7.2e-16
C11_202 341 329 7.2e-16
R11_21 344 343 0.001
C11_211 344 329 2.4e-16
C11_212 343 329 2.4e-16
R11_22 345 344 0.001
C11_221 345 329 2.4e-16
C11_222 344 329 2.4e-16
R11_23 340 345 0.3
C11_231 340 329 4.44e-15
C11_232 345 329 4.44e-15
R11_24 338 340 0.1
C11_241 338 329 2.28e-15
C11_242 340 329 2.28e-15
R11_25 337 338 0.001
C11_251 337 329 1.32e-15
C11_252 338 329 1.32e-15
R11_26 334 337 0.1
C11_261 334 329 1.56e-15
C11_262 337 329 1.56e-15
R11_27 335 334 0.001
C11_271 335 329 7.2e-16
C11_272 334 329 7.2e-16
R11_28 336 335 0.001
C11_281 336 329 2.4e-16
C11_282 335 329 2.4e-16
R11_29 332 336 0.001
C11_291 332 329 3.6e-16
C11_292 336 329 3.6e-16
R11_30 333 332 0.1
C11_301 333 329 2.28e-15
C11_302 332 329 2.28e-15
R11_31 328 333 0.001
C11_311 328 329 7.2e-16
C11_312 333 329 7.2e-16
R11_32 327 328 0.001
C11_321 327 329 3.9e-16
C11_322 328 329 3.9e-16
R11_33 325 327 0.1
C11_331 325 329 7.605e-15
C11_332 327 329 7.605e-15
R11_34 326 325 0.001
C11_341 326 329 3.705e-15
C11_342 325 329 3.705e-15
R11_35 320 326 0.001
C11_351 320 329 2.145e-15
C11_352 326 329 2.145e-15
R11_36 321 320 0.001
C11_361 321 329 2.535e-15
C11_362 320 329 2.535e-15
R11_37 322 321 0.001
C11_371 322 329 1.17e-15
C11_372 321 329 1.17e-15
R11_38 313 312 0.001
C11_381 313 329 3.705e-15
C11_382 312 329 3.705e-15
R11_39 312 329 0.001
C11_391 312 329 1.2e-15
C11_392 329 329 1.2e-15
R11_40 313 329 0.001
C11_401 313 329 1.08e-15
C11_402 329 329 1.08e-15
R11_41 315 313 0.001
C11_411 315 329 1.56e-15
C11_412 313 329 1.56e-15
R11_42 323 322 0.001
C11_421 323 329 3.9e-16
C11_422 322 329 3.9e-16
R11_43 324 323 0.001
C11_431 324 329 3.9e-16
C11_432 323 329 3.9e-16
R11_44 319 324 0.1
C11_441 319 329 7.215e-15
C11_442 324 329 7.215e-15
R11_45 318 319 0.001
C11_451 318 329 3.705e-15
C11_452 319 329 3.705e-15
R11_46 312 316 0.001
C11_461 312 329 5.85e-16
C11_462 316 329 5.85e-16
R11_47 317 318 0.001
C11_471 317 329 2.145e-15
C11_472 318 329 2.145e-15
R11_48 311 317 0.001
C11_481 311 329 2.535e-15
C11_482 317 329 2.535e-15
R11_49 314 311 0.001
C11_491 314 329 1.17e-15
C11_492 311 329 1.17e-15
R11_50 316 314 0.001
C11_501 316 329 3.9e-16
C11_502 314 329 3.9e-16
R10_1 361 360 0.001
R10_2 360 362 0.9
C10_21 360 329 1.0925e-15
C10_22 362 329 1.0925e-15
R10_3 358 360 1.5
C10_31 358 329 1.7825e-15
C10_32 360 329 1.7825e-15
R10_4 361 363 500
C10_41 361 329 1.5e-15
C10_42 363 329 1.5e-15
R10_5 359 361 550
C10_51 359 329 1.65e-15
C10_52 361 329 1.65e-15
R8_1 369 379 0.001
R8_2 369 378 0.001
R8_3 381 380 0.001
R8_4 383 384 0.001
R8_5 375 374 400
C8_51 375 329 1.275e-15
C8_52 374 329 1.275e-15
R8_6 376 375 50
C8_61 376 329 1.5e-16
C8_62 375 329 1.5e-16
R8_7 377 376 50
C8_71 377 329 2.25e-16
C8_72 376 329 2.25e-16
R8_8 372 377 700
C8_81 372 329 2.175e-15
C8_82 377 329 2.175e-15
R8_9 373 372 50
C8_91 373 329 1.5e-16
C8_92 372 329 1.5e-16
R8_10 371 373 300
C8_101 371 329 9.75e-16
C8_102 373 329 9.75e-16
R8_11 371 382 1200
C8_111 371 329 3.6e-15
C8_112 382 329 3.6e-15
R8_12 381 382 200
C8_121 381 329 6e-16
C8_122 382 329 6e-16
R8_13 380 384 0.5
C8_131 380 329 1.4e-15
C8_132 384 329 1.4e-15
R8_14 379 380 0.5
C8_141 379 329 1.4e-15
C8_142 380 329 1.4e-15
R8_15 378 379 0.2
C8_151 378 329 7e-16
C8_152 379 329 7e-16
R8_16 370 378 0.2
C8_161 370 329 7.7e-16
C8_162 378 329 7.7e-16
R7_1 390 389 0.001
R7_2 389 391 0.9
C7_21 389 329 1.0925e-15
C7_22 391 329 1.0925e-15
R7_3 387 389 1.5
C7_31 387 329 1.7825e-15
C7_32 389 329 1.7825e-15
R7_4 390 392 500
C7_41 390 329 1.5e-15
C7_42 392 329 1.5e-15
R7_5 388 390 550
C7_51 388 329 1.65e-15
C7_52 390 329 1.65e-15
R6_1 395 396 0.001
R6_2 408 407 0.001
R6_3 411 412 0.001
R6_4 410 409 0.001
R6_5 415 416 0.001
R6_6 401 402 0.001
R6_7 425 424 0.001
R6_8 424 426 0.001
R6_9 426 423 550
C6_91 426 329 1.65e-15
C6_92 423 329 1.65e-15
R6_10 420 426 500
C6_101 420 329 1.5e-15
C6_102 426 329 1.5e-15
R6_11 424 427 1.5
C6_111 424 329 1.7825e-15
C6_112 427 329 1.7825e-15
R6_12 421 424 0.9
C6_121 421 329 1.0925e-15
C6_122 424 329 1.0925e-15
R6_13 422 425 0.3
C6_131 422 329 1.44e-15
C6_132 425 329 1.44e-15
R6_14 402 403 0.1
C6_141 402 329 1.725e-16
C6_142 403 329 1.725e-16
R6_15 405 402 0.2
C6_151 405 329 2.875e-16
C6_152 402 329 2.875e-16
R6_16 417 416 0.1
C6_161 417 329 1.725e-16
C6_162 416 329 1.725e-16
R6_17 419 422 2.3
C6_171 419 329 1.104e-14
C6_172 422 329 1.104e-14
R6_18 418 417 0.1
C6_181 418 329 1.15e-16
C6_182 417 329 1.15e-16
R6_19 409 418 0.9
C6_191 409 329 1.0925e-15
C6_192 418 329 1.0925e-15
R6_20 404 409 1
C6_201 404 329 1.2075e-15
C6_202 409 329 1.2075e-15
R6_21 403 404 0.1
C6_211 403 329 1.15e-16
C6_212 404 329 1.15e-16
R6_22 410 419 0.8
C6_221 410 329 3.84e-15
C6_222 419 329 3.84e-15
R6_23 406 410 0.15
C6_231 406 329 8.4e-16
C6_232 410 329 8.4e-16
R6_24 397 406 1.1
C6_241 397 329 5.4e-15
C6_242 406 329 5.4e-15
R6_25 397 408 0.15
C6_251 397 329 8.4e-16
C6_252 408 329 8.4e-16
R6_26 413 412 0.1
C6_261 413 329 1.725e-16
C6_262 412 329 1.725e-16
R6_27 414 413 0.1
C6_271 414 329 1.15e-16
C6_272 413 329 1.15e-16
R6_28 407 414 0.9
C6_281 407 329 1.0925e-15
C6_282 414 329 1.0925e-15
R6_29 398 407 1
C6_291 398 329 1.2075e-15
C6_292 407 329 1.2075e-15
R6_30 399 398 0.1
C6_301 399 329 1.15e-16
C6_302 398 329 1.15e-16
R6_31 396 399 0.1
C6_311 396 329 1.725e-16
C6_312 399 329 1.725e-16
R6_32 400 396 0.2
C6_321 400 329 2.875e-16
C6_322 396 329 2.875e-16
R4_1 440 439 0.001
R4_2 438 437 0.001
R4_3 479 477 0.001
R4_4 473 472 0.001
R4_5 475 474 0.001
R4_6 442 441 0.001
R4_7 474 476 0.001
R4_8 441 443 0.001
R4_9 450 455 200
C4_91 450 329 6.75e-16
C4_92 455 329 6.75e-16
R4_10 464 471 200
C4_101 464 329 6.75e-16
C4_102 471 329 6.75e-16
R4_11 456 457 50
C4_111 456 329 2.25e-16
C4_112 457 329 2.25e-16
R4_12 455 456 50
C4_121 455 329 1.5e-16
C4_122 456 329 1.5e-16
R4_13 465 464 50
C4_131 465 329 1.5e-16
C4_132 464 329 1.5e-16
R4_14 466 465 50
C4_141 466 329 2.25e-16
C4_142 465 329 2.25e-16
R4_15 453 457 700
C4_151 453 329 2.175e-15
C4_152 457 329 2.175e-15
R4_16 462 466 700
C4_161 462 329 2.175e-15
C4_162 466 329 2.175e-15
R4_17 454 453 50
C4_171 454 329 1.5e-16
C4_172 453 329 1.5e-16
R4_18 451 454 300
C4_181 451 329 9.75e-16
C4_182 454 329 9.75e-16
R4_19 463 462 50
C4_191 463 329 1.5e-16
C4_192 462 329 1.5e-16
R4_20 460 463 300
C4_201 460 329 9.75e-16
C4_202 463 329 9.75e-16
R4_21 452 451 100
C4_211 452 329 3e-16
C4_212 451 329 3e-16
R4_22 460 461 100
C4_221 460 329 3e-16
C4_222 461 329 3e-16
R4_23 447 452 400
C4_231 447 329 1.2e-15
C4_232 452 329 1.2e-15
R4_24 459 461 400
C4_241 459 329 1.2e-15
C4_242 461 329 1.2e-15
R4_25 443 447 450
C4_251 443 329 1.35e-15
C4_252 447 329 1.35e-15
R4_26 435 443 700
C4_261 435 329 2.1e-15
C4_262 443 329 2.1e-15
R4_27 476 480 700
C4_271 476 329 2.1e-15
C4_272 480 329 2.1e-15
R4_28 459 476 450
C4_281 459 329 1.35e-15
C4_282 476 329 1.35e-15
R4_29 473 478 700
C4_291 473 329 2.1e-15
C4_292 478 329 2.1e-15
R4_30 458 473 450
C4_301 458 329 1.35e-15
C4_302 473 329 1.35e-15
R4_31 441 448 0.5
C4_311 441 329 1.47e-15
C4_312 448 329 1.47e-15
R4_32 436 441 1
C4_321 436 329 2.87e-15
C4_322 441 329 2.87e-15
R4_33 474 482 1
C4_331 474 329 2.87e-15
C4_332 482 329 2.87e-15
R4_34 469 474 0.5
C4_341 469 329 1.47e-15
C4_342 474 329 1.47e-15
R4_35 442 449 0.1
C4_351 442 329 6e-16
C4_352 449 329 6e-16
R4_36 470 475 0.1
C4_361 470 329 6e-16
C4_362 475 329 6e-16
R4_37 477 481 0.6
C4_371 477 329 1.75e-15
C4_372 481 329 1.75e-15
R4_38 472 477 0.4
C4_381 472 329 1.12e-15
C4_382 477 329 1.12e-15
R4_39 467 472 0.5
C4_391 467 329 1.47e-15
C4_392 472 329 1.47e-15
R4_40 445 449 1.5
C4_401 445 329 7.2e-15
C4_402 449 329 7.2e-15
R4_41 468 470 1.5
C4_411 468 329 7.2e-15
C4_412 470 329 7.2e-15
R4_42 468 479 0.3
C4_421 468 329 1.56e-15
C4_422 479 329 1.56e-15
R4_43 445 468 0.75
C4_431 445 329 3.6e-15
C4_432 468 329 3.6e-15
R4_44 438 445 0.3
C4_441 438 329 1.56e-15
C4_442 445 329 1.56e-15
R4_45 439 446 0.5
C4_451 439 329 1.47e-15
C4_452 446 329 1.47e-15
R4_46 437 439 0.4
C4_461 437 329 1.12e-15
C4_462 439 329 1.12e-15
R4_47 434 437 0.6
C4_471 434 329 1.75e-15
C4_472 437 329 1.75e-15
R4_48 440 444 450
C4_481 440 329 1.35e-15
C4_482 444 329 1.35e-15
R4_49 433 440 700
C4_491 433 329 2.1e-15
C4_492 440 329 2.1e-15
R3_1 485 495 0.001
R3_2 485 494 0.001
R3_3 497 496 0.001
R3_4 499 500 0.001
R3_5 491 490 400
C3_51 491 329 1.275e-15
C3_52 490 329 1.275e-15
R3_6 492 491 50
C3_61 492 329 1.5e-16
C3_62 491 329 1.5e-16
R3_7 493 492 50
C3_71 493 329 2.25e-16
C3_72 492 329 2.25e-16
R3_8 488 493 700
C3_81 488 329 2.175e-15
C3_82 493 329 2.175e-15
R3_9 489 488 50
C3_91 489 329 1.5e-16
C3_92 488 329 1.5e-16
R3_10 487 489 300
C3_101 487 329 9.75e-16
C3_102 489 329 9.75e-16
R3_11 487 498 1200
C3_111 487 329 3.6e-15
C3_112 498 329 3.6e-15
R3_12 497 498 200
C3_121 497 329 6e-16
C3_122 498 329 6e-16
R3_13 496 500 0.5
C3_131 496 329 1.4e-15
C3_132 500 329 1.4e-15
R3_14 495 496 0.5
C3_141 495 329 1.4e-15
C3_142 496 329 1.4e-15
R3_15 494 495 0.2
C3_151 494 329 7e-16
C3_152 495 329 7e-16
R3_16 486 494 0.2
C3_161 486 329 7.7e-16
C3_162 494 329 7.7e-16
R2_1 509 510 0.001
R2_2 514 515 0.001
R2_3 504 506 0.001
R2_4 517 518 0.001
R2_5 524 525 0.001
R2_6 525 526 0.3
C2_61 525 329 4.92e-15
C2_62 526 329 4.92e-15
R2_7 523 525 0.1
C2_71 523 329 2.28e-15
C2_72 525 329 2.28e-15
R2_8 522 523 0.001
C2_81 522 329 1.32e-15
C2_82 523 329 1.32e-15
R2_9 518 522 0.1
C2_91 518 329 1.56e-15
C2_92 522 329 1.56e-15
R2_10 519 518 0.001
C2_101 519 329 7.2e-16
C2_102 518 329 7.2e-16
R2_11 507 505 0.001
C2_111 507 329 7.2e-16
C2_112 505 329 7.2e-16
R2_12 507 503 0.001
C2_121 507 329 4.8e-16
C2_122 503 329 4.8e-16
R2_13 506 503 0.001
C2_131 506 329 1.08e-15
C2_132 503 329 1.08e-15
R2_14 508 506 0.001
C2_141 508 329 9.6e-16
C2_142 506 329 9.6e-16
R2_15 520 519 0.001
C2_151 520 329 2.4e-16
C2_152 519 329 2.4e-16
R2_16 521 520 0.001
C2_161 521 329 2.4e-16
C2_162 520 329 2.4e-16
R2_17 515 521 0.3
C2_171 515 329 4.44e-15
C2_172 521 329 4.44e-15
R2_18 516 515 0.1
C2_181 516 329 2.28e-15
C2_182 515 329 2.28e-15
R2_19 505 512 0.001
C2_191 505 329 3.6e-16
C2_192 512 329 3.6e-16
R2_20 511 516 0.001
C2_201 511 329 1.32e-15
C2_202 516 329 1.32e-15
R2_21 510 511 0.1
C2_211 510 329 1.56e-15
C2_212 511 329 1.56e-15
R2_22 513 510 0.001
C2_221 513 329 7.2e-16
C2_222 510 329 7.2e-16
R2_23 512 513 0.001
C2_231 512 329 2.4e-16
C2_232 513 329 2.4e-16
R1_1 529 534 0.001
R1_2 529 533 0.001
R1_3 542 543 0.001
R1_4 535 534 0.001
R1_5 538 537 0.001
R1_6 537 539 0.001
R1_7 541 549 200
C1_71 541 329 6.75e-16
C1_72 549 329 6.75e-16
R1_8 550 551 50
C1_81 550 329 2.25e-16
C1_82 551 329 2.25e-16
R1_9 549 550 50
C1_91 549 329 1.5e-16
C1_92 550 329 1.5e-16
R1_10 547 551 700
C1_101 547 329 2.175e-15
C1_102 551 329 2.175e-15
R1_11 548 547 50
C1_111 548 329 1.5e-16
C1_112 547 329 1.5e-16
R1_12 545 548 300
C1_121 545 329 9.75e-16
C1_122 548 329 9.75e-16
R1_13 546 545 100
C1_131 546 329 3e-16
C1_132 545 329 3e-16
R1_14 540 546 400
C1_141 540 329 1.2e-15
C1_142 546 329 1.2e-15
R1_15 539 540 450
C1_151 539 329 1.35e-15
C1_152 540 329 1.35e-15
R1_16 532 539 700
C1_161 532 329 2.1e-15
C1_162 539 329 2.1e-15
R1_17 537 544 0.5
C1_171 537 329 1.47e-15
C1_172 544 329 1.47e-15
R1_18 531 537 1
C1_181 531 329 2.87e-15
C1_182 537 329 2.87e-15
R1_19 536 538 0.2
C1_191 536 329 9.6e-16
C1_192 538 329 9.6e-16
R1_20 535 536 0.25
C1_201 535 329 1.2e-15
C1_202 536 329 1.2e-15
R1_21 534 543 0.9
C1_211 534 329 2.66e-15
C1_212 543 329 2.66e-15
R1_22 533 534 0.3
C1_221 533 329 8.4e-16
C1_222 534 329 8.4e-16
R1_23 530 533 0.2
C1_231 530 329 7.7e-16
C1_232 533 329 7.7e-16
.ends mux4inv

