.include mux.spi

x1 10 11 12 20 30 40 mux

v1 11 30 sine(0.9 0.9 0.25G 0 0 0)
v2 10 30 pulse(0 1.8 0ns 1ns 1ns 1ps 2ns)
v3 12 30 pulse(0 1.8 0ns 1ps 1ps 8ns 16ns)
v4 20 30 1.8V
v5 30 0 0V DC

.tran 0.001ns 16ns

.model tp pmos level=54
.model tn nmos level=54

.end 
