module inv(input logic [3:0] a, output logic [3:0] saida);
     assign saida=~a;
endmodule