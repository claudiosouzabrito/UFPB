* Spice description of mux4
* Spice driver version 348321288
* Date ( dd/mm/yyyy hh:mm:ss ):  6/08/2019 at 14:41:28

* INTERF d0 d1 d2 d3 s0 s1 vdd vdd2 vss y 


.subckt mux4 209 166 280 273 387 105 43 404 266 58 
* NET 1 = mux3.tiristor2.inversor_1.vdd
* NET 9 = mux3.tiristor1.inversor_1.vdd
* NET 23 = mux1.tiristor2.inversor_1.vdd
* NET 43 = vdd
* NET 58 = y
* NET 74 = mux3.tiristor2.inversor_1.vss
* NET 105 = s1
* NET 118 = mux3.inversor.inversor_1.nq
* NET 152 = mux3.inversor.inversor_1.vss
* NET 166 = d1
* NET 209 = d0
* NET 214 = mux2.tiristor2.inversor_1.vss
* NET 222 = mux1.inversor.inversor_1.nq
* NET 266 = vss
* NET 273 = d3
* NET 280 = d2
* NET 321 = mux2.tiristor2.inversor_1.vdd
* NET 387 = s0
* NET 404 = vdd2
* NET 416 = mux2.tiristor1.inversor_1.nq
Mtr_00036 109 141 1 404 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00035 315 142 64 404 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00034 139 107 10 404 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00033 193 108 60 404 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00032 136 104 9 404 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00031 9 104 136 404 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00030 335 419 321 404 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00029 271 422 291 404 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00028 424 332 406 404 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00027 278 334 285 404 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00026 416 329 401 404 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00025 401 329 416 404 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00024 392 245 23 404 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00023 167 246 191 404 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00022 243 390 32 404 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00021 210 391 189 404 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00020 240 388 31 404 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00019 31 388 240 404 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00018 74 125 85 266 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00017 312 88 51 266 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00016 157 84 120 266 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00015 179 123 46 266 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00014 152 81 118 266 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00013 152 81 118 266 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00012 214 444 360 266 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00011 274 356 306 266 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00010 257 359 442 266 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00009 281 438 301 266 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00008 256 344 440 266 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00007 256 344 440 266 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00006 219 229 371 266 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00005 164 374 175 266 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00004 268 365 224 266 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00003 207 227 171 266 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00002 267 364 222 266 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00001 267 364 222 266 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
R22_1 1 2 0.001
R22_2 5 6 0.001
C22_21 5 266 6e-16
C22_22 6 266 6e-16
R22_3 4 5 0.001
C22_31 4 266 7.2e-16
C22_32 5 266 7.2e-16
R22_4 2 4 0.1
C22_41 2 266 1.44e-15
C22_42 4 266 1.44e-15
R22_5 3 2 0.001
C22_51 3 266 1.08e-15
C22_52 2 266 1.08e-15
R21_1 10 17 0.001
R21_2 9 11 0.001
R21_3 14 15 0.001
C21_31 14 266 3.6e-16
C21_32 15 266 3.6e-16
R21_4 13 14 0.001
C21_41 13 266 7.2e-16
C21_42 14 266 7.2e-16
R21_5 11 13 0.1
C21_51 11 266 1.56e-15
C21_52 13 266 1.56e-15
R21_6 12 11 0.001
C21_61 12 266 9.6e-16
C21_62 11 266 9.6e-16
R21_7 18 20 0.001
C21_71 18 266 6e-16
C21_72 20 266 6e-16
R21_8 19 18 0.001
C21_81 19 266 7.2e-16
C21_82 18 266 7.2e-16
R21_9 17 19 0.1
C21_91 17 266 1.44e-15
C21_92 19 266 1.44e-15
R21_10 16 17 0.001
C21_101 16 266 8.4e-16
C21_102 17 266 8.4e-16
R21_11 15 16 0.001
C21_111 15 266 2.4e-16
C21_112 16 266 2.4e-16
R20_1 23 24 0.001
R20_2 27 28 0.001
C20_21 27 266 6e-16
C20_22 28 266 6e-16
R20_3 26 27 0.001
C20_31 26 266 7.2e-16
C20_32 27 266 7.2e-16
R20_4 24 26 0.1
C20_41 24 266 1.44e-15
C20_42 26 266 1.44e-15
R20_5 25 24 0.001
C20_51 25 266 1.08e-15
C20_52 24 266 1.08e-15
R19_1 32 39 0.001
R19_2 31 33 0.001
R19_3 36 37 0.001
C19_31 36 266 3.6e-16
C19_32 37 266 3.6e-16
R19_4 35 36 0.001
C19_41 35 266 7.2e-16
C19_42 36 266 7.2e-16
R19_5 35 43 0.001
C19_51 35 266 4.8e-16
C19_52 43 266 4.8e-16
R19_6 33 43 0.001
C19_61 33 266 1.08e-15
C19_62 43 266 1.08e-15
R19_7 34 33 0.001
C19_71 34 266 9.6e-16
C19_72 33 266 9.6e-16
R19_8 40 42 0.001
C19_81 40 266 6e-16
C19_82 42 266 6e-16
R19_9 41 40 0.001
C19_91 41 266 7.2e-16
C19_92 40 266 7.2e-16
R19_10 39 41 0.1
C19_101 39 266 1.44e-15
C19_102 41 266 1.44e-15
R19_11 38 39 0.001
C19_111 38 266 8.4e-16
C19_112 39 266 8.4e-16
R19_12 37 38 0.001
C19_121 37 266 2.4e-16
C19_122 38 266 2.4e-16
R18_1 46 47 0.001
R18_2 57 56 0.001
R18_3 60 68 0.001
R18_4 59 58 0.001
R18_5 64 70 0.001
R18_6 51 52 0.001
R18_7 52 53 0.1
C18_71 52 266 1.725e-16
C18_72 53 266 1.725e-16
R18_8 55 52 0.2
C18_81 55 266 2.875e-16
C18_82 52 266 2.875e-16
R18_9 70 71 0.2
C18_91 70 266 2.875e-16
C18_92 71 266 2.875e-16
R18_10 65 70 0.1
C18_101 65 266 1.725e-16
C18_102 70 266 1.725e-16
R18_11 66 65 0.1
C18_111 66 266 1.15e-16
C18_112 65 266 1.15e-16
R18_12 58 66 1
C18_121 58 266 1.2075e-15
C18_122 66 266 1.2075e-15
R18_13 54 58 0.9
C18_131 54 266 1.0925e-15
C18_132 58 266 1.0925e-15
R18_14 53 54 0.1
C18_141 53 266 1.15e-16
C18_142 54 266 1.15e-16
R18_15 59 67 0.15
C18_151 59 266 8.4e-16
C18_152 67 266 8.4e-16
R18_16 61 67 0.75
C18_161 61 266 3.6e-15
C18_162 67 266 3.6e-15
R18_17 57 61 0.15
C18_171 57 266 8.4e-16
C18_172 61 266 8.4e-16
R18_18 68 69 0.2
C18_181 68 266 2.875e-16
C18_182 69 266 2.875e-16
R18_19 62 68 0.1
C18_191 62 266 1.725e-16
C18_192 68 266 1.725e-16
R18_20 63 62 0.1
C18_201 63 266 1.15e-16
C18_202 62 266 1.15e-16
R18_21 56 63 1
C18_211 56 266 1.2075e-15
C18_212 63 266 1.2075e-15
R18_22 48 56 0.9
C18_221 48 266 1.0925e-15
C18_222 56 266 1.0925e-15
R18_23 49 48 0.1
C18_231 49 266 1.15e-16
C18_232 48 266 1.15e-16
R18_24 47 49 0.1
C18_241 47 266 1.725e-16
C18_242 49 266 1.725e-16
R18_25 50 47 0.2
C18_251 50 266 2.875e-16
C18_252 47 266 2.875e-16
R17_1 74 75 0.001
R17_2 77 78 0.001
C17_21 77 266 6e-16
C17_22 78 266 6e-16
R17_3 75 77 0.1
C17_31 75 266 2.16e-15
C17_32 77 266 2.16e-15
R17_4 76 75 0.001
C17_41 76 266 1.08e-15
C17_42 75 266 1.08e-15
R16_1 93 92 0.001
R16_2 106 105 0.001
R16_3 96 95 0.001
R16_4 95 97 0.001
R16_5 100 99 0.001
R16_6 99 101 0.001
R16_7 109 111 0.001
R16_8 109 110 0.001
R16_9 85 86 0.001
R16_10 89 88 250
C16_101 89 266 7.5e-16
C16_102 88 266 7.5e-16
R16_11 87 89 350
C16_111 87 266 1.05e-15
C16_112 89 266 1.05e-15
R16_12 87 102 650
C16_121 87 266 1.95e-15
C16_122 102 266 1.95e-15
R16_13 101 102 200
C16_131 101 266 6e-16
C16_132 102 266 6e-16
R16_14 114 108 750
C16_141 114 266 2.25e-15
C16_142 108 266 2.25e-15
R16_15 107 114 450
C16_151 107 266 1.425e-15
C16_152 114 266 1.425e-15
R16_16 111 115 0.2
C16_161 111 266 7.7e-16
C16_162 115 266 7.7e-16
R16_17 110 111 0.2
C16_171 110 266 7e-16
C16_172 111 266 7e-16
R16_18 99 110 0.5
C16_181 99 266 1.4e-15
C16_182 110 266 1.4e-15
R16_19 86 99 0.5
C16_191 86 266 1.4e-15
C16_192 99 266 1.4e-15
R16_20 97 107 600
C16_201 97 266 1.875e-15
C16_202 107 266 1.875e-15
R16_21 84 97 500
C16_211 84 266 1.5e-15
C16_212 97 266 1.5e-15
R16_22 103 100 0.1
C16_221 103 266 4.8e-16
C16_222 100 266 4.8e-16
R16_23 91 103 0.05
C16_231 91 266 2.4e-16
C16_232 103 266 2.4e-16
R16_24 90 91 0.85
C16_241 90 266 4.2e-15
C16_242 91 266 4.2e-15
R16_25 95 113 1
C16_251 95 266 2.87e-15
C16_252 113 266 2.87e-15
R16_26 83 95 0.5
C16_261 83 266 1.47e-15
C16_262 95 266 1.47e-15
R16_27 98 96 0.05
C16_271 98 266 3.6e-16
C16_272 96 266 3.6e-16
R16_28 90 98 0.05
C16_281 90 266 3.6e-16
C16_282 98 266 3.6e-16
R16_29 94 96 0.35
C16_291 94 266 1.8e-15
C16_292 96 266 1.8e-15
R16_30 94 106 0.2
C16_301 94 266 9.6e-16
C16_302 106 266 9.6e-16
R16_31 105 112 0.6
C16_311 105 266 1.75e-15
C16_312 112 266 1.75e-15
R16_32 92 105 0.4
C16_321 92 266 1.12e-15
C16_322 105 266 1.12e-15
R16_33 82 92 0.5
C16_331 82 266 1.47e-15
C16_332 92 266 1.47e-15
R16_34 93 104 700
C16_341 93 266 2.1e-15
C16_342 104 266 2.1e-15
R16_35 81 93 450
C16_351 81 266 1.35e-15
C16_352 93 266 1.35e-15
R15_1 118 119 0.001
R15_2 136 144 0.001
R15_3 136 137 0.001
R15_4 138 137 0.001
R15_5 128 127 0.001
R15_6 127 129 0.001
R15_7 139 145 0.001
R15_8 139 143 0.001
R15_9 120 121 0.001
R15_10 133 132 0.001
R15_11 132 134 0.001
R15_12 148 142 750
C15_121 148 266 2.25e-15
C15_122 142 266 2.25e-15
R15_13 141 148 450
C15_131 141 266 1.425e-15
C15_132 148 266 1.425e-15
R15_14 134 141 600
C15_141 134 266 1.875e-15
C15_142 141 266 1.875e-15
R15_15 125 134 500
C15_151 125 266 1.5e-15
C15_152 134 266 1.5e-15
R15_16 124 123 250
C15_161 124 266 7.5e-16
C15_162 123 266 7.5e-16
R15_17 122 124 350
C15_171 122 266 1.05e-15
C15_172 124 266 1.05e-15
R15_18 132 149 1
C15_181 132 266 2.87e-15
C15_182 149 266 2.87e-15
R15_19 126 132 0.5
C15_191 126 266 1.47e-15
C15_192 132 266 1.47e-15
R15_20 122 130 650
C15_201 122 266 1.95e-15
C15_202 130 266 1.95e-15
R15_21 129 130 200
C15_211 129 266 6e-16
C15_212 130 266 6e-16
R15_22 135 133 0.05
C15_221 135 266 3.6e-16
C15_222 133 266 3.6e-16
R15_23 131 135 0.6
C15_231 131 266 3e-15
C15_232 135 266 3e-15
R15_24 145 147 0.2
C15_241 145 266 7.7e-16
C15_242 147 266 7.7e-16
R15_25 143 145 0.2
C15_251 143 266 7e-16
C15_252 145 266 7e-16
R15_26 127 143 0.5
C15_261 127 266 1.4e-15
C15_262 143 266 1.4e-15
R15_27 121 127 0.5
C15_271 121 266 1.4e-15
C15_272 127 266 1.4e-15
R15_28 131 128 0.05
C15_281 131 266 3.6e-16
C15_282 128 266 3.6e-16
R15_29 128 140 0.2
C15_291 128 266 9.6e-16
C15_292 140 266 9.6e-16
R15_30 138 140 0.35
C15_301 138 266 1.8e-15
C15_302 140 266 1.8e-15
R15_31 144 146 0.2
C15_311 144 266 7.7e-16
C15_312 146 266 7.7e-16
R15_32 137 144 0.3
C15_321 137 266 8.4e-16
C15_322 144 266 8.4e-16
R15_33 119 137 0.9
C15_331 119 266 2.66e-15
C15_332 137 266 2.66e-15
R14_1 152 153 0.001
R14_2 157 158 0.001
R14_3 160 161 0.001
C14_31 160 266 6e-16
C14_32 161 266 6e-16
R14_4 158 160 0.1
C14_41 158 266 2.16e-15
C14_42 160 266 2.16e-15
R14_5 159 158 0.001
C14_51 159 266 8.4e-16
C14_52 158 266 8.4e-16
R14_6 156 159 0.001
C14_61 156 266 2.4e-16
C14_62 159 266 2.4e-16
R14_7 155 156 0.001
C14_71 155 266 3.6e-16
C14_72 156 266 3.6e-16
R14_8 153 155 0.1
C14_81 153 266 2.28e-15
C14_82 155 266 2.28e-15
R14_9 154 153 0.001
C14_91 154 266 9.6e-16
C14_92 153 266 9.6e-16
R13_1 164 165 0.001
R13_2 167 168 0.001
R13_3 166 168 1.3
C13_31 166 266 1.495e-15
C13_32 168 266 1.495e-15
R13_4 165 166 1.2
C13_41 165 266 1.38e-15
C13_42 166 266 1.38e-15
R12_1 171 172 0.001
R12_2 184 183 0.001
R12_3 189 194 0.001
R12_4 186 185 0.001
R12_5 188 187 0.001
R12_6 191 197 0.001
R12_7 175 176 0.001
R12_8 193 200 0.001
R12_9 179 180 0.001
R12_10 187 200 1.3
C12_101 187 266 1.495e-15
C12_102 200 266 1.495e-15
R12_11 180 187 1.2
C12_111 180 266 1.38e-15
C12_112 187 266 1.38e-15
R12_12 176 177 0.1
C12_121 176 266 1.725e-16
C12_122 177 266 1.725e-16
R12_13 178 176 0.2
C12_131 178 266 2.875e-16
C12_132 176 266 2.875e-16
R12_14 197 203 0.2
C12_141 197 266 2.875e-16
C12_142 203 266 2.875e-16
R12_15 198 197 0.1
C12_151 198 266 1.725e-16
C12_152 197 266 1.725e-16
R12_16 188 204 0.35
C12_161 188 266 1.68e-15
C12_162 204 266 1.68e-15
R12_17 199 198 0.1
C12_171 199 266 1.15e-16
C12_172 198 266 1.15e-16
R12_18 185 199 1
C12_181 185 266 1.2075e-15
C12_182 199 266 1.2075e-15
R12_19 182 185 0.9
C12_191 182 266 1.0925e-15
C12_192 185 266 1.0925e-15
R12_20 177 182 0.1
C12_201 177 266 1.15e-16
C12_202 182 266 1.15e-16
R12_21 202 204 0.95
C12_211 202 266 4.68e-15
C12_212 204 266 4.68e-15
R12_22 192 202 0.15
C12_221 192 266 8.4e-16
C12_222 202 266 8.4e-16
R12_23 186 192 0.15
C12_231 186 266 8.4e-16
C12_232 192 266 8.4e-16
R12_24 190 192 0.75
C12_241 190 266 3.6e-15
C12_242 192 266 3.6e-15
R12_25 184 190 0.15
C12_251 184 266 8.4e-16
C12_252 190 266 8.4e-16
R12_26 194 201 0.2
C12_261 194 266 2.875e-16
C12_262 201 266 2.875e-16
R12_27 195 194 0.1
C12_271 195 266 1.725e-16
C12_272 194 266 1.725e-16
R12_28 196 195 0.1
C12_281 196 266 1.15e-16
C12_282 195 266 1.15e-16
R12_29 183 196 1
C12_291 183 266 1.2075e-15
C12_292 196 266 1.2075e-15
R12_30 181 183 0.9
C12_301 181 266 1.0925e-15
C12_302 183 266 1.0925e-15
R12_31 173 181 0.1
C12_311 173 266 1.15e-16
C12_312 181 266 1.15e-16
R12_32 172 173 0.1
C12_321 172 266 1.725e-16
C12_322 173 266 1.725e-16
R12_33 174 172 0.2
C12_331 174 266 2.875e-16
C12_332 172 266 2.875e-16
R11_1 207 208 0.001
R11_2 210 211 0.001
R11_3 209 211 1.3
C11_31 209 266 1.495e-15
C11_32 211 266 1.495e-15
R11_4 208 209 1.2
C11_41 208 266 1.38e-15
C11_42 209 266 1.38e-15
R10_1 214 215 0.001
R10_2 219 215 0.001
R10_3 217 218 0.001
C10_31 217 266 9.75e-16
C10_32 218 266 9.75e-16
R10_4 215 217 0.001
C10_41 215 266 3.51e-15
C10_42 217 266 3.51e-15
R10_5 216 215 0.001
C10_51 216 266 1.755e-15
C10_52 215 266 1.755e-15
R9_1 222 223 0.001
R9_2 240 248 0.001
R9_3 240 241 0.001
R9_4 242 241 0.001
R9_5 232 231 0.001
R9_6 231 233 0.001
R9_7 243 249 0.001
R9_8 243 247 0.001
R9_9 224 225 0.001
R9_10 237 236 0.001
R9_11 236 238 0.001
R9_12 252 246 750
C9_121 252 266 2.25e-15
C9_122 246 266 2.25e-15
R9_13 245 252 450
C9_131 245 266 1.425e-15
C9_132 252 266 1.425e-15
R9_14 238 245 600
C9_141 238 266 1.875e-15
C9_142 245 266 1.875e-15
R9_15 229 238 500
C9_151 229 266 1.5e-15
C9_152 238 266 1.5e-15
R9_16 228 227 250
C9_161 228 266 7.5e-16
C9_162 227 266 7.5e-16
R9_17 226 228 350
C9_171 226 266 1.05e-15
C9_172 228 266 1.05e-15
R9_18 236 253 1
C9_181 236 266 2.87e-15
C9_182 253 266 2.87e-15
R9_19 230 236 0.5
C9_191 230 266 1.47e-15
C9_192 236 266 1.47e-15
R9_20 226 234 650
C9_201 226 266 1.95e-15
C9_202 234 266 1.95e-15
R9_21 233 234 200
C9_211 233 266 6e-16
C9_212 234 266 6e-16
R9_22 239 237 0.05
C9_221 239 266 3.6e-16
C9_222 237 266 3.6e-16
R9_23 235 239 0.6
C9_231 235 266 3e-15
C9_232 239 266 3e-15
R9_24 249 251 0.2
C9_241 249 266 7.7e-16
C9_242 251 266 7.7e-16
R9_25 247 249 0.2
C9_251 247 266 7e-16
C9_252 249 266 7e-16
R9_26 231 247 0.5
C9_261 231 266 1.4e-15
C9_262 247 266 1.4e-15
R9_27 225 231 0.5
C9_271 225 266 1.4e-15
C9_272 231 266 1.4e-15
R9_28 235 232 0.05
C9_281 235 266 3.6e-16
C9_282 232 266 3.6e-16
R9_29 232 244 0.2
C9_291 232 266 9.6e-16
C9_292 244 266 9.6e-16
R9_30 242 244 0.35
C9_301 242 266 1.8e-15
C9_302 244 266 1.8e-15
R9_31 248 250 0.2
C9_311 248 266 7.7e-16
C9_312 250 266 7.7e-16
R9_32 241 248 0.3
C9_321 241 266 8.4e-16
C9_322 248 266 8.4e-16
R9_33 223 241 0.9
C9_331 223 266 2.66e-15
C9_332 241 266 2.66e-15
R8_1 256 258 0.001
R8_2 257 262 0.001
R8_3 268 262 0.001
R8_4 267 258 0.001
R8_5 258 260 0.001
C8_51 258 266 3.705e-15
C8_52 260 266 3.705e-15
R8_6 264 265 0.001
C8_61 264 266 9.75e-16
C8_62 265 266 9.75e-16
R8_7 262 264 0.001
C8_71 262 266 3.51e-15
C8_72 264 266 3.51e-15
R8_8 263 262 0.001
C8_81 263 266 1.365e-15
C8_82 262 266 1.365e-15
R8_9 261 263 0.001
C8_91 261 266 3.9e-16
C8_92 263 266 3.9e-16
R8_10 260 261 0.001
C8_101 260 266 5.85e-16
C8_102 261 266 5.85e-16
R8_11 260 266 0.001
C8_111 260 266 1.2e-15
C8_112 266 266 1.2e-15
R8_12 258 266 0.001
C8_121 258 266 1.08e-15
C8_122 266 266 1.08e-15
R8_13 259 258 0.001
C8_131 259 266 1.56e-15
C8_132 258 266 1.56e-15
R7_1 271 272 0.001
R7_2 274 275 0.001
R7_3 273 275 1.2
C7_31 273 266 1.38e-15
C7_32 275 266 1.38e-15
R7_4 272 273 1.3
C7_41 272 266 1.495e-15
C7_42 273 266 1.495e-15
R6_1 278 279 0.001
R6_2 281 282 0.001
R6_3 280 282 1.2
C6_31 280 266 1.38e-15
C6_32 282 266 1.38e-15
R6_4 279 280 1.3
C6_41 279 266 1.495e-15
C6_42 280 266 1.495e-15
R5_1 285 286 0.001
R5_2 298 297 0.001
R5_3 301 302 0.001
R5_4 300 299 0.001
R5_5 306 307 0.001
R5_6 291 292 0.001
R5_7 317 316 0.001
R5_8 315 318 0.001
R5_9 312 313 0.001
R5_10 316 318 1.3
C5_101 316 266 1.495e-15
C5_102 318 266 1.495e-15
R5_11 313 316 1.2
C5_111 313 266 1.38e-15
C5_112 316 266 1.38e-15
R5_12 314 317 0.25
C5_121 314 266 1.32e-15
C5_122 317 266 1.32e-15
R5_13 292 293 0.1
C5_131 292 266 1.725e-16
C5_132 293 266 1.725e-16
R5_14 295 292 0.2
C5_141 295 266 2.875e-16
C5_142 292 266 2.875e-16
R5_15 307 309 0.2
C5_151 307 266 2.875e-16
C5_152 309 266 2.875e-16
R5_16 308 307 0.1
C5_161 308 266 1.725e-16
C5_162 307 266 1.725e-16
R5_17 311 314 1.7
C5_171 311 266 8.28e-15
C5_172 314 266 8.28e-15
R5_18 310 308 0.1
C5_181 310 266 1.15e-16
C5_182 308 266 1.15e-16
R5_19 299 310 0.9
C5_191 299 266 1.0925e-15
C5_192 310 266 1.0925e-15
R5_20 294 299 1
C5_201 294 266 1.2075e-15
C5_202 299 266 1.2075e-15
R5_21 293 294 0.1
C5_211 293 266 1.15e-16
C5_212 294 266 1.15e-16
R5_22 300 311 0.8
C5_221 300 266 3.96e-15
C5_222 311 266 3.96e-15
R5_23 296 300 0.15
C5_231 296 266 8.4e-16
C5_232 300 266 8.4e-16
R5_24 287 296 0.75
C5_241 287 266 3.6e-15
C5_242 296 266 3.6e-15
R5_25 287 298 0.15
C5_251 287 266 8.4e-16
C5_252 298 266 8.4e-16
R5_26 302 304 0.2
C5_261 302 266 2.875e-16
C5_262 304 266 2.875e-16
R5_27 303 302 0.1
C5_271 303 266 1.725e-16
C5_272 302 266 1.725e-16
R5_28 305 303 0.1
C5_281 305 266 1.15e-16
C5_282 303 266 1.15e-16
R5_29 297 305 0.9
C5_291 297 266 1.0925e-15
C5_292 305 266 1.0925e-15
R5_30 288 297 1
C5_301 288 266 1.2075e-15
C5_302 297 266 1.2075e-15
R5_31 289 288 0.1
C5_311 289 266 1.15e-16
C5_312 288 266 1.15e-16
R5_32 286 289 0.1
C5_321 286 266 1.725e-16
C5_322 289 266 1.725e-16
R5_33 290 286 0.2
C5_331 290 266 2.875e-16
C5_332 286 266 2.875e-16
R4_1 321 322 0.001
R4_2 325 326 0.001
C4_21 325 266 6e-16
C4_22 326 266 6e-16
R4_3 324 325 0.001
C4_31 324 266 7.2e-16
C4_32 325 266 7.2e-16
R4_4 322 324 0.1
C4_41 322 266 1.44e-15
C4_42 324 266 1.44e-15
R4_5 323 322 0.001
C4_51 323 266 1.08e-15
C4_52 322 266 1.08e-15
R3_1 342 347 0.001
R3_2 347 348 0.001
R3_3 339 338 0.001
R3_4 389 387 0.001
R3_5 352 351 0.001
R3_6 379 378 0.001
R3_7 351 343 0.001
R3_8 341 345 0.001
R3_9 376 375 0.001
R3_10 378 380 0.001
R3_11 360 361 0.001
R3_12 335 340 0.001
R3_13 335 336 0.001
R3_14 383 382 0.001
R3_15 382 384 0.001
R3_16 392 393 0.001
R3_17 392 394 0.001
R3_18 371 372 0.001
R3_19 367 374 250
C3_191 367 266 7.5e-16
C3_192 374 266 7.5e-16
R3_20 366 367 350
C3_201 366 266 1.05e-15
C3_202 367 266 1.05e-15
R3_21 366 386 650
C3_211 366 266 1.95e-15
C3_212 386 266 1.95e-15
R3_22 384 386 200
C3_221 384 266 6e-16
C3_222 386 266 6e-16
R3_23 397 391 750
C3_231 397 266 2.25e-15
C3_232 391 266 2.25e-15
R3_24 356 363 250
C3_241 356 266 7.5e-16
C3_242 363 266 7.5e-16
R3_25 390 397 450
C3_251 390 266 1.425e-15
C3_252 397 266 1.425e-15
R3_26 362 363 350
C3_261 362 266 1.05e-15
C3_262 363 266 1.05e-15
R3_27 393 398 0.2
C3_271 393 266 7.7e-16
C3_272 398 266 7.7e-16
R3_28 394 393 0.2
C3_281 394 266 7e-16
C3_282 393 266 7e-16
R3_29 382 394 0.5
C3_291 382 266 1.4e-15
C3_292 394 266 1.4e-15
R3_30 372 382 0.5
C3_301 372 266 1.4e-15
C3_302 382 266 1.4e-15
R3_31 380 390 600
C3_311 380 266 1.875e-15
C3_312 390 266 1.875e-15
R3_32 365 380 500
C3_321 365 266 1.5e-15
C3_322 380 266 1.5e-15
R3_33 355 362 650
C3_331 355 266 1.95e-15
C3_332 362 266 1.95e-15
R3_34 376 388 700
C3_341 376 266 2.1e-15
C3_342 388 266 2.1e-15
R3_35 364 376 450
C3_351 364 266 1.35e-15
C3_352 376 266 1.35e-15
R3_36 341 344 450
C3_361 341 266 1.35e-15
C3_362 344 266 1.35e-15
R3_37 329 341 700
C3_371 329 266 2.1e-15
C3_372 341 266 2.1e-15
R3_38 343 355 200
C3_381 343 266 6e-16
C3_382 355 266 6e-16
R3_39 385 383 0.1
C3_391 385 266 4.8e-16
C3_392 383 266 4.8e-16
R3_40 373 385 0.05
C3_401 373 266 2.4e-16
C3_402 385 266 2.4e-16
R3_41 369 373 0.85
C3_411 369 266 4.2e-15
C3_412 373 266 4.2e-15
R3_42 378 396 1
C3_421 378 266 2.87e-15
C3_422 396 266 2.87e-15
R3_43 370 378 0.5
C3_431 370 266 1.47e-15
C3_432 378 266 1.47e-15
R3_44 351 361 0.5
C3_441 351 266 1.4e-15
C3_442 361 266 1.4e-15
R3_45 340 351 0.5
C3_451 340 266 1.4e-15
C3_452 351 266 1.4e-15
R3_46 336 340 0.2
C3_461 336 266 7e-16
C3_462 340 266 7e-16
R3_47 337 336 0.2
C3_471 337 266 7.7e-16
C3_472 336 266 7.7e-16
R3_48 381 379 0.05
C3_481 381 266 3.6e-16
C3_482 379 266 3.6e-16
R3_49 369 381 0.05
C3_491 369 266 3.6e-16
C3_492 381 266 3.6e-16
R3_50 387 395 0.6
C3_501 387 266 1.75e-15
C3_502 395 266 1.75e-15
R3_51 375 387 0.4
C3_511 375 266 1.12e-15
C3_512 387 266 1.12e-15
R3_52 368 375 0.5
C3_521 368 266 1.47e-15
C3_522 375 266 1.47e-15
R3_53 345 357 0.5
C3_531 345 266 1.47e-15
C3_532 357 266 1.47e-15
R3_54 338 345 0.4
C3_541 338 266 1.12e-15
C3_542 345 266 1.12e-15
R3_55 330 338 0.6
C3_551 330 266 1.75e-15
C3_552 338 266 1.75e-15
R3_56 377 379 0.35
C3_561 377 266 1.8e-15
C3_562 379 266 1.8e-15
R3_57 352 353 0.1
C3_571 352 266 4.8e-16
C3_572 353 266 4.8e-16
R3_58 353 354 0.05
C3_581 353 266 2.4e-16
C3_582 354 266 2.4e-16
R3_59 377 389 0.2
C3_591 377 266 9.6e-16
C3_592 389 266 9.6e-16
R3_60 346 377 1
C3_601 346 266 4.8e-15
C3_602 377 266 4.8e-15
R3_61 339 346 0.2
C3_611 339 266 9.6e-16
C3_612 346 266 9.6e-16
R3_62 349 354 0.85
C3_621 349 266 4.2e-15
C3_622 354 266 4.2e-15
R3_63 346 348 0.35
C3_631 346 266 1.8e-15
C3_632 348 266 1.8e-15
R3_64 350 349 0.05
C3_641 350 266 3.6e-16
C3_642 349 266 3.6e-16
R3_65 348 350 0.05
C3_651 348 266 3.6e-16
C3_652 350 266 3.6e-16
R3_66 333 334 750
C3_661 333 266 2.25e-15
C3_662 334 266 2.25e-15
R3_67 347 358 0.5
C3_671 347 266 1.47e-15
C3_672 358 266 1.47e-15
R3_68 331 347 1
C3_681 331 266 2.87e-15
C3_682 347 266 2.87e-15
R3_69 333 332 450
C3_691 333 266 1.425e-15
C3_692 332 266 1.425e-15
R3_70 342 359 500
C3_701 342 266 1.5e-15
C3_702 359 266 1.5e-15
R3_71 332 342 600
C3_711 332 266 1.875e-15
C3_712 342 266 1.875e-15
R2_1 406 410 0.001
R2_2 401 402 0.001
R2_3 407 408 0.001
C2_31 407 266 3.6e-16
C2_32 408 266 3.6e-16
R2_4 405 407 0.001
C2_41 405 266 7.2e-16
C2_42 407 266 7.2e-16
R2_5 405 404 0.001
C2_51 405 266 4.8e-16
C2_52 404 266 4.8e-16
R2_6 402 404 0.001
C2_61 402 266 1.08e-15
C2_62 404 266 1.08e-15
R2_7 403 402 0.001
C2_71 403 266 9.6e-16
C2_72 402 266 9.6e-16
R2_8 411 413 0.001
C2_81 411 266 6e-16
C2_82 413 266 6e-16
R2_9 412 411 0.001
C2_91 412 266 7.2e-16
C2_92 411 266 7.2e-16
R2_10 410 412 0.1
C2_101 410 266 1.44e-15
C2_102 412 266 1.44e-15
R2_11 409 410 0.001
C2_111 409 266 8.4e-16
C2_112 410 266 8.4e-16
R2_12 408 409 0.001
C2_121 408 266 2.4e-16
C2_122 409 266 2.4e-16
R1_1 424 428 0.001
R1_2 424 425 0.001
R1_3 431 430 0.001
R1_4 442 443 0.001
R1_5 432 430 0.001
R1_6 427 426 0.001
R1_7 435 434 0.001
R1_8 434 436 0.001
R1_9 440 441 0.001
R1_10 416 426 0.001
R1_11 416 423 0.001
R1_12 420 422 750
C1_121 420 266 2.25e-15
C1_122 422 266 2.25e-15
R1_13 420 419 450
C1_131 420 266 1.425e-15
C1_132 419 266 1.425e-15
R1_14 436 444 500
C1_141 436 266 1.5e-15
C1_142 444 266 1.5e-15
R1_15 419 436 600
C1_151 419 266 1.875e-15
C1_152 436 266 1.875e-15
R1_16 434 447 0.5
C1_161 434 266 1.47e-15
C1_162 447 266 1.47e-15
R1_17 421 434 1
C1_171 421 266 2.87e-15
C1_172 434 266 2.87e-15
R1_18 426 441 0.9
C1_181 426 266 2.66e-15
C1_182 441 266 2.66e-15
R1_19 423 426 0.3
C1_191 423 266 8.4e-16
C1_192 426 266 8.4e-16
R1_20 417 423 0.2
C1_201 417 266 7.7e-16
C1_202 423 266 7.7e-16
R1_21 438 446 250
C1_211 438 266 7.5e-16
C1_212 446 266 7.5e-16
R1_22 435 439 0.05
C1_221 435 266 3.6e-16
C1_222 439 266 3.6e-16
R1_23 445 446 350
C1_231 445 266 1.05e-15
C1_232 446 266 1.05e-15
R1_24 427 429 0.35
C1_241 427 266 1.8e-15
C1_242 429 266 1.8e-15
R1_25 437 439 0.6
C1_251 437 266 3e-15
C1_252 439 266 3e-15
R1_26 433 445 650
C1_261 433 266 1.95e-15
C1_262 445 266 1.95e-15
R1_27 429 432 0.2
C1_271 429 266 9.6e-16
C1_272 432 266 9.6e-16
R1_28 432 437 0.05
C1_281 432 266 3.6e-16
C1_282 437 266 3.6e-16
R1_29 431 433 200
C1_291 431 266 6e-16
C1_292 433 266 6e-16
R1_30 430 443 0.5
C1_301 430 266 1.4e-15
C1_302 443 266 1.4e-15
R1_31 428 430 0.5
C1_311 428 266 1.4e-15
C1_312 430 266 1.4e-15
R1_32 425 428 0.2
C1_321 425 266 7e-16
C1_322 428 266 7e-16
R1_33 418 425 0.2
C1_331 418 266 7.7e-16
C1_332 425 266 7.7e-16
.ends mux4

