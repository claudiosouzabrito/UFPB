.subckt c1 1 2
C1 1 2 1u
.ends c1
