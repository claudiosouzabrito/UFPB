* Spice description of biel8
* Spice driver version 1140717064
* Date ( dd/mm/yyyy hh:mm:ss ):  9/07/2019 at 12:41:50

* INTERF a vdd vss y y2 y3 


.subckt biel8 27 50 82 58 15 2 
* NET 2 = y3
* NET 15 = y2
* NET 27 = a
* NET 50 = vdd
* NET 58 = y
* NET 82 = vss
Mtr_00006 38 22 5 50 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00005 37 65 20 50 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00004 36 33 63 50 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00003 1 13 77 82 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00002 10 56 74 82 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00001 53 31 70 82 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
R6_1 1 3 0.001
R6_2 5 6 0.001
R6_3 6 7 0.4
C6_31 6 82 1.33e-15
C6_32 7 82 1.33e-15
R6_4 2 6 0.6
C6_41 2 82 1.82e-15
C6_42 6 82 1.82e-15
R6_5 3 2 0.2
C6_51 3 82 7e-16
C6_52 2 82 7e-16
R6_6 4 3 0.1
C6_61 4 82 4.9e-16
C6_62 3 82 4.9e-16
R5_1 10 11 0.001
R5_2 20 21 0.001
R5_3 18 17 0.001
R5_4 18 22 700
C5_41 18 82 2.1e-15
C5_42 22 82 2.1e-15
R5_5 13 18 300
C5_51 13 82 9e-16
C5_52 18 82 9e-16
R5_6 19 24 0.8
C5_61 19 82 2.45e-15
C5_62 24 82 2.45e-15
R5_7 17 19 0.1
C5_71 17 82 4.2e-16
C5_72 19 82 4.2e-16
R5_8 14 17 0.5
C5_81 14 82 1.47e-15
C5_82 17 82 1.47e-15
R5_9 16 19 1.5
C5_91 16 82 1.725e-15
C5_92 19 82 1.725e-15
R5_10 21 23 0.4
C5_101 21 82 1.33e-15
C5_102 23 82 1.33e-15
R5_11 16 21 0.4
C5_111 16 82 1.12e-15
C5_112 21 82 1.12e-15
R5_12 15 16 0.2
C5_121 15 82 7e-16
C5_122 16 82 7e-16
R5_13 11 15 0.2
C5_131 11 82 7e-16
C5_132 15 82 7e-16
R5_14 12 11 0.1
C5_141 12 82 4.9e-16
C5_142 11 82 4.9e-16
R4_1 29 28 0.001
R4_2 28 32 1
C4_21 28 82 2.87e-15
C4_22 32 82 2.87e-15
R4_3 27 28 0.1
C4_31 27 82 4.2e-16
C4_32 28 82 4.2e-16
R4_4 30 27 0.3
C4_41 30 82 1.05e-15
C4_42 27 82 1.05e-15
R4_5 29 33 700
C4_51 29 82 2.1e-15
C4_52 33 82 2.1e-15
R4_6 31 29 300
C4_61 31 82 9e-16
C4_62 29 82 9e-16
R3_1 36 39 0.001
R3_2 37 42 0.001
R3_3 38 45 0.001
R3_4 48 49 0.001
C3_41 48 82 6e-16
C3_42 49 82 6e-16
R3_5 50 48 0.1
C3_51 50 82 1.68e-15
C3_52 48 82 1.68e-15
R3_6 45 50 0.001
C3_61 45 82 7.2e-16
C3_62 50 82 7.2e-16
R3_7 46 45 0.001
C3_71 46 82 3.6e-16
C3_72 45 82 3.6e-16
R3_8 47 46 0.001
C3_81 47 82 2.4e-16
C3_82 46 82 2.4e-16
R3_9 44 47 0.1
C3_91 44 82 1.8e-15
C3_92 47 82 1.8e-15
R3_10 42 44 0.1
C3_101 42 82 2.4e-15
C3_102 44 82 2.4e-15
R3_11 43 42 0.001
C3_111 43 82 6e-16
C3_112 42 82 6e-16
R3_12 40 43 0.2
C3_121 40 82 3e-15
C3_122 43 82 3e-15
R3_13 39 40 0.1
C3_131 39 82 2.4e-15
C3_132 40 82 2.4e-15
R3_14 41 39 0.001
C3_141 41 82 6e-16
C3_142 39 82 6e-16
R2_1 53 54 0.001
R2_2 63 64 0.001
R2_3 61 60 0.001
R2_4 61 65 700
C2_41 61 82 2.1e-15
C2_42 65 82 2.1e-15
R2_5 56 61 300
C2_51 56 82 9e-16
C2_52 61 82 9e-16
R2_6 62 67 0.8
C2_61 62 82 2.45e-15
C2_62 67 82 2.45e-15
R2_7 60 62 0.1
C2_71 60 82 4.2e-16
C2_72 62 82 4.2e-16
R2_8 57 60 0.5
C2_81 57 82 1.47e-15
C2_82 60 82 1.47e-15
R2_9 59 62 2
C2_91 59 82 2.3e-15
C2_92 62 82 2.3e-15
R2_10 64 66 0.4
C2_101 64 82 1.33e-15
C2_102 66 82 1.33e-15
R2_11 59 64 0.4
C2_111 59 82 1.12e-15
C2_112 64 82 1.12e-15
R2_12 58 59 0.2
C2_121 58 82 7e-16
C2_122 59 82 7e-16
R2_13 54 58 0.2
C2_131 54 82 7e-16
C2_132 58 82 7e-16
R2_14 55 54 0.1
C2_141 55 82 4.9e-16
C2_142 54 82 4.9e-16
R1_1 70 71 0.001
R1_2 74 75 0.001
R1_3 77 79 0.001
R1_4 83 84 0.001
C1_41 83 82 6e-16
C1_42 84 82 6e-16
R1_5 83 82 0.1
C1_51 83 82 1.44e-15
C1_52 82 82 1.44e-15
R1_6 79 82 0.001
C1_61 79 82 7.2e-16
C1_62 82 82 7.2e-16
R1_7 80 79 0.001
C1_71 80 82 6e-16
C1_72 79 82 6e-16
R1_8 81 80 0.001
C1_81 81 82 2.4e-16
C1_82 80 82 2.4e-16
R1_9 78 81 0.1
C1_91 78 82 1.8e-15
C1_92 81 82 1.8e-15
R1_10 75 78 0.1
C1_101 75 82 2.16e-15
C1_102 78 82 2.16e-15
R1_11 76 75 0.001
C1_111 76 82 8.4e-16
C1_112 75 82 8.4e-16
R1_12 72 76 0.2
C1_121 72 82 3e-15
C1_122 76 82 3e-15
R1_13 71 72 0.1
C1_131 71 82 2.16e-15
C1_132 72 82 2.16e-15
R1_14 73 71 0.001
C1_141 73 82 8.4e-16
C1_142 71 82 8.4e-16
.ends biel8

