* Spice description of transmissiongate2
* Spice driver version -1435929080
* Date ( dd/mm/yyyy hh:mm:ss ): 29/07/2019 at 13:41:25

* INTERF a s vdd vss y 


.subckt transmissiongate2 34 3 16 56 25 
* NET 3 = s
* NET 16 = vdd
* NET 25 = y
* NET 34 = a
* NET 39 = inversor_1.nq
* NET 56 = vss
Mtr_00006 47 5 10 16 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00005 10 5 47 16 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00004 35 6 24 16 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00003 53 1 39 56 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00002 53 1 39 56 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00001 32 42 19 56 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
R6_1 4 3 0.001
R6_2 3 7 1
C6_21 3 56 2.87e-15
C6_22 7 56 2.87e-15
R6_3 2 3 0.5
C6_31 2 56 1.47e-15
C6_32 3 56 1.47e-15
R6_4 5 6 750
C6_41 5 56 2.25e-15
C6_42 6 56 2.25e-15
R6_5 4 5 700
C6_51 4 56 2.1375e-15
C6_52 5 56 2.1375e-15
R6_6 1 4 450
C6_61 1 56 1.35e-15
C6_62 4 56 1.35e-15
R5_1 10 11 0.001
R5_2 14 15 0.001
C5_21 14 56 6e-16
C5_22 15 56 6e-16
R5_3 13 14 0.001
C5_31 13 56 7.2e-16
C5_32 14 56 7.2e-16
R5_4 13 16 0.001
C5_41 13 56 4.8e-16
C5_42 16 56 4.8e-16
R5_5 11 16 0.001
C5_51 11 56 1.08e-15
C5_52 16 56 1.08e-15
R5_6 12 11 0.001
C5_61 12 56 9.6e-16
C5_62 11 56 9.6e-16
R4_1 19 20 0.001
R4_2 24 26 0.001
R4_3 26 28 0.2
C4_31 26 56 2.875e-16
C4_32 28 56 2.875e-16
R4_4 27 26 0.1
C4_41 27 56 1.725e-16
C4_42 26 56 1.725e-16
R4_5 29 27 0.1
C4_51 29 56 1.15e-16
C4_52 27 56 1.15e-16
R4_6 25 29 1
C4_61 25 56 1.2075e-15
C4_62 29 56 1.2075e-15
R4_7 21 25 0.9
C4_71 21 56 1.0925e-15
C4_72 25 56 1.0925e-15
R4_8 22 21 0.1
C4_81 22 56 1.15e-16
C4_82 21 56 1.15e-16
R4_9 20 22 0.1
C4_91 20 56 1.725e-16
C4_92 22 56 1.725e-16
R4_10 23 20 0.2
C4_101 23 56 2.875e-16
C4_102 20 56 2.875e-16
R3_1 32 33 0.001
R3_2 35 36 0.001
R3_3 34 36 1.3
C3_31 34 56 1.495e-15
C3_32 36 56 1.495e-15
R3_4 33 34 1.2
C3_41 33 56 1.38e-15
C3_42 34 56 1.38e-15
R2_1 39 40 0.001
R2_2 47 49 0.001
R2_3 47 48 0.001
R2_4 45 44 0.001
R2_5 43 42 250
C2_51 43 56 7.5e-16
C2_52 42 56 7.5e-16
R2_6 41 43 350
C2_61 41 56 1.05e-15
C2_62 43 56 1.05e-15
R2_7 41 46 650
C2_71 41 56 1.95e-15
C2_72 46 56 1.95e-15
R2_8 45 46 200
C2_81 45 56 6e-16
C2_82 46 56 6e-16
R2_9 49 50 0.2
C2_91 49 56 7.7e-16
C2_92 50 56 7.7e-16
R2_10 48 49 0.2
C2_101 48 56 7e-16
C2_102 49 56 7e-16
R2_11 44 48 0.5
C2_111 44 56 1.4e-15
C2_112 48 56 1.4e-15
R2_12 40 44 0.5
C2_121 40 56 1.4e-15
C2_122 44 56 1.4e-15
R1_1 53 54 0.001
R1_2 57 58 0.001
C1_21 57 56 6e-16
C1_22 58 56 6e-16
R1_3 57 56 0.001
C1_31 57 56 1.2e-15
C1_32 56 56 1.2e-15
R1_4 54 56 0.001
C1_41 54 56 1.08e-15
C1_42 56 56 1.08e-15
R1_5 55 54 0.001
C1_51 55 56 9.6e-16
C1_52 54 56 9.6e-16
.ends transmissiongate2

