module inv(input logic a, output logic saida);
     assign saida=~a;
endmodule