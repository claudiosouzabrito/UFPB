
.include nand2.spi
.model tp pmos level=54
.model tn nmos level=54

x1 10 11 20 30 40 nand2

v1 10 30 0V DC

v2 11 30 1.8v DC

v3 20 30 1.8v DC
v4 30 0 0v

.dc v1 0 +1.8 0.001
.end
