* Spice description of flipflop
* Spice driver version -1620904440
* Date ( dd/mm/yyyy hh:mm:ss ): 15/08/2019 at 15:51:30

* INTERF clk d q vdd vss 


.subckt flipflop 167 116 23 214 273 
* NET 23 = q
* NET 29 = latch2.inv1.nq
* NET 46 = latch2.mux.i0
* NET 93 = latch1.inv1.nq
* NET 116 = d
* NET 119 = latch1.mux.q
* NET 167 = clk
* NET 183 = latch1.mux.i0
* NET 214 = vdd
* NET 253 = inv.nq
* NET 273 = vss
Mtr_00034 262 166 199 214 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00033 191 99 203 214 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00032 100 133 202 214 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00031 200 154 134 214 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00030 7 114 200 214 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00029 316 265 208 214 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00028 10 266 156 214 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00027 156 318 7 214 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00026 208 188 10 214 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00025 54 35 207 214 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00024 36 21 206 214 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00023 204 73 19 214 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00022 4 136 204 214 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00021 87 178 210 214 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00020 1 177 75 214 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00019 75 89 4 214 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00018 210 51 1 214 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00017 300 161 253 273 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00016 302 96 184 273 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00015 301 120 93 273 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00014 297 110 146 273 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00013 146 256 149 273 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00012 296 255 309 273 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00011 149 311 250 273 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00010 250 183 296 273 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00009 119 150 297 273 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00008 304 32 47 273 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00007 303 16 29 273 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00006 299 121 65 273 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00005 65 163 68 273 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00004 298 164 80 273 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00003 68 82 62 273 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00002 62 46 298 273 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00001 13 69 299 273 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
R19_1 13 14 0.001
R19_2 19 22 0.001
R19_3 19 23 0.001
R19_4 24 23 0.001
R19_5 19 20 0.001
R19_6 26 25 0.001
R19_7 18 17 0.001
R19_8 18 21 600
C19_81 18 273 1.875e-15
C19_82 21 273 1.875e-15
R19_9 16 18 500
C19_91 16 273 1.5e-15
C19_92 18 273 1.5e-15
R19_10 17 25 1
C19_101 17 273 2.8e-15
C19_102 25 273 2.8e-15
R19_11 15 17 0.5
C19_111 15 273 1.47e-15
C19_112 17 273 1.47e-15
R19_12 24 26 0.25
C19_121 24 273 1.2e-15
C19_122 26 273 1.2e-15
R19_13 22 23 0.2
C19_131 22 273 7e-16
C19_132 23 273 7e-16
R19_14 20 22 0.2
C19_141 20 273 7e-16
C19_142 22 273 7e-16
R19_15 14 20 1
C19_151 14 273 2.8e-15
C19_152 20 273 2.8e-15
R18_1 29 30 0.001
R18_2 36 38 0.001
R18_3 39 38 0.001
R18_4 36 37 0.001
R18_5 41 40 0.001
R18_6 34 33 0.001
R18_7 34 35 600
C18_71 34 273 1.875e-15
C18_72 35 273 1.875e-15
R18_8 32 34 500
C18_81 32 273 1.5e-15
C18_82 34 273 1.5e-15
R18_9 40 43 0.2
C18_91 40 273 7.7e-16
C18_92 43 273 7.7e-16
R18_10 33 40 0.7
C18_101 33 273 2.1e-15
C18_102 40 273 2.1e-15
R18_11 31 33 0.5
C18_111 31 273 1.47e-15
C18_112 33 273 1.47e-15
R18_12 39 41 0.25
C18_121 39 273 1.2e-15
C18_122 41 273 1.2e-15
R18_13 38 42 0.2
C18_131 38 273 7.7e-16
C18_132 42 273 7.7e-16
R18_14 37 38 0.2
C18_141 37 273 7e-16
C18_142 38 273 7e-16
R18_15 30 37 1
C18_151 30 273 2.8e-15
C18_152 37 273 2.8e-15
R17_1 50 49 0.001
R17_2 51 52 0.001
R17_3 53 52 0.001
R17_4 56 55 0.001
R17_5 55 54 0.001
R17_6 54 57 0.001
R17_7 47 48 0.001
R17_8 57 59 0.2
C17_81 57 273 7.7e-16
C17_82 59 273 7.7e-16
R17_9 55 57 0.2
C17_91 55 273 7e-16
C17_92 57 273 7e-16
R17_10 48 55 1
C17_101 48 273 2.8e-15
C17_102 55 273 2.8e-15
R17_11 53 56 1.5
C17_111 53 273 7.2e-15
C17_112 56 273 7.2e-15
R17_12 52 58 0.5
C17_121 52 273 1.47e-15
C17_122 58 273 1.47e-15
R17_13 49 52 0.7
C17_131 49 273 2.1e-15
C17_132 52 273 2.1e-15
R17_14 46 50 500
C17_141 46 273 1.5e-15
C17_142 50 273 1.5e-15
R14_1 68 70 0.001
R14_2 75 76 0.001
R14_3 75 77 0.001
R14_4 72 71 0.001
R14_5 74 73 700
C14_51 74 273 2.175e-15
C14_52 73 273 2.175e-15
R14_6 69 74 750
C14_61 69 273 2.325e-15
C14_62 74 273 2.325e-15
R14_7 72 74 900
C14_71 72 273 2.7e-15
C14_72 74 273 2.7e-15
R14_8 76 77 0.5
C14_81 76 273 5.75e-16
C14_82 77 273 5.75e-16
R14_9 71 76 1.1
C14_91 71 273 1.265e-15
C14_92 76 273 1.265e-15
R14_10 70 71 0.9
C14_101 70 273 1.035e-15
C14_102 71 273 1.035e-15
R13_1 80 81 0.001
R13_2 82 83 0.001
R13_3 87 90 0.001
R13_4 87 88 0.001
R13_5 86 85 0.001
R13_6 86 89 500
C13_61 86 273 1.575e-15
C13_62 89 273 1.575e-15
R13_7 84 85 1.7
C13_71 84 273 1.955e-15
C13_72 85 273 1.955e-15
R13_8 88 90 0.5
C13_81 88 273 5.75e-16
C13_82 90 273 5.75e-16
R13_9 81 88 2.5
C13_91 81 273 2.875e-15
C13_92 88 273 2.875e-15
R13_10 83 84 0.9
C13_101 83 273 1.035e-15
C13_102 84 273 1.035e-15
R13_11 81 83 1.3
C13_111 81 273 1.495e-15
C13_112 83 273 1.495e-15
R12_1 93 94 0.001
R12_2 100 102 0.001
R12_3 103 102 0.001
R12_4 100 101 0.001
R12_5 105 104 0.001
R12_6 98 97 0.001
R12_7 98 99 600
C12_71 98 273 1.875e-15
C12_72 99 273 1.875e-15
R12_8 96 98 500
C12_81 96 273 1.5e-15
C12_82 98 273 1.5e-15
R12_9 104 107 0.2
C12_91 104 273 7.7e-16
C12_92 107 273 7.7e-16
R12_10 97 104 0.7
C12_101 97 273 2.1e-15
C12_102 104 273 2.1e-15
R12_11 95 97 0.5
C12_111 95 273 1.47e-15
C12_112 97 273 1.47e-15
R12_12 103 105 0.25
C12_121 103 273 1.2e-15
C12_122 105 273 1.2e-15
R12_13 102 106 0.2
C12_131 102 273 7.7e-16
C12_132 106 273 7.7e-16
R12_14 101 102 0.2
C12_141 101 273 7e-16
C12_142 102 273 7e-16
R12_15 94 101 1
C12_151 94 273 2.8e-15
C12_152 101 273 2.8e-15
R11_1 111 112 0.001
R11_2 114 115 0.001
R11_3 115 116 0.5
C11_31 115 273 1.4e-15
C11_32 116 273 1.4e-15
R11_4 112 115 0.7
C11_41 112 273 2.1e-15
C11_42 115 273 2.1e-15
R11_5 113 112 0.2
C11_51 113 273 7.7e-16
C11_52 112 273 7.7e-16
R11_6 110 111 500
C11_61 110 273 1.5e-15
C11_62 111 273 1.5e-15
R10_1 119 122 0.001
R10_2 134 138 0.001
R10_3 134 139 0.001
R10_4 140 139 0.001
R10_5 134 135 0.001
R10_6 128 127 0.001
R10_7 142 141 0.001
R10_8 132 131 0.001
R10_9 130 129 0.001
R10_10 125 124 0.001
R10_11 136 137 0.001
R10_12 121 125 500
C10_121 121 273 1.5e-15
C10_122 125 273 1.5e-15
R10_13 130 133 600
C10_131 130 273 1.875e-15
C10_132 133 273 1.875e-15
R10_14 120 130 500
C10_141 120 273 1.5e-15
C10_142 130 273 1.5e-15
R10_15 137 143 0.5
C10_151 137 273 1.47e-15
C10_152 143 273 1.47e-15
R10_16 131 137 0.5
C10_161 131 273 1.4e-15
C10_162 137 273 1.4e-15
R10_17 124 131 0.2
C10_171 124 273 7e-16
C10_172 131 273 7e-16
R10_18 126 124 0.2
C10_181 126 273 7.7e-16
C10_182 124 273 7.7e-16
R10_19 129 141 1
C10_191 129 273 2.8e-15
C10_192 141 273 2.8e-15
R10_20 123 129 0.5
C10_201 123 273 1.47e-15
C10_202 129 273 1.47e-15
R10_21 128 132 1.6
C10_211 128 273 7.8e-15
C10_212 132 273 7.8e-15
R10_22 140 142 0.25
C10_221 140 273 1.2e-15
C10_222 142 273 1.2e-15
R10_23 138 139 0.2
C10_231 138 273 7e-16
C10_232 139 273 7e-16
R10_24 135 138 0.2
C10_241 135 273 7e-16
C10_242 138 273 7e-16
R10_25 127 135 0.5
C10_251 127 273 1.4e-15
C10_252 135 273 1.4e-15
R10_26 122 127 0.5
C10_261 122 273 1.4e-15
C10_262 127 273 1.4e-15
R8_1 149 151 0.001
R8_2 156 157 0.001
R8_3 156 158 0.001
R8_4 153 152 0.001
R8_5 155 154 700
C8_51 155 273 2.175e-15
C8_52 154 273 2.175e-15
R8_6 150 155 750
C8_61 150 273 2.325e-15
C8_62 155 273 2.325e-15
R8_7 153 155 900
C8_71 153 273 2.7e-15
C8_72 155 273 2.7e-15
R8_8 157 158 0.5
C8_81 157 273 5.75e-16
C8_82 158 273 5.75e-16
R8_9 152 157 1.1
C8_91 152 273 1.265e-15
C8_92 157 273 1.265e-15
R8_10 151 152 0.9
C8_101 151 273 1.035e-15
C8_102 152 273 1.035e-15
R7_1 169 168 0.001
R7_2 170 167 0.001
R7_3 172 171 0.001
R7_4 174 173 0.001
R7_5 175 178 850
C7_51 175 273 2.625e-15
C7_52 178 273 2.625e-15
R7_6 164 175 750
C7_61 164 273 2.25e-15
C7_62 175 273 2.25e-15
R7_7 163 176 750
C7_71 163 273 2.25e-15
C7_72 176 273 2.25e-15
R7_8 174 177 850
C7_81 174 273 2.625e-15
C7_82 177 273 2.625e-15
R7_9 174 176 450
C7_91 174 273 1.35e-15
C7_92 176 273 1.35e-15
R7_10 175 174 450
C7_101 175 273 1.35e-15
C7_102 174 273 1.35e-15
R7_11 171 180 0.7
C7_111 171 273 2.17e-15
C7_112 180 273 2.17e-15
R7_12 173 171 0.2
C7_121 173 273 7e-16
C7_122 171 273 7e-16
R7_13 165 173 0.2
C7_131 165 273 7.7e-16
C7_132 173 273 7.7e-16
R7_14 170 172 2.5
C7_141 170 273 1.2e-14
C7_142 172 273 1.2e-14
R7_15 167 179 0.7
C7_151 167 273 2.17e-15
C7_152 179 273 2.17e-15
R7_16 168 167 0.2
C7_161 168 273 7e-16
C7_162 167 273 7e-16
R7_17 162 168 0.5
C7_171 162 273 1.47e-15
C7_172 168 273 1.47e-15
R7_18 169 166 600
C7_181 169 273 1.875e-15
C7_182 166 273 1.875e-15
R7_19 161 169 500
C7_191 161 273 1.5e-15
C7_192 169 273 1.5e-15
R6_1 187 186 0.001
R6_2 188 189 0.001
R6_3 190 189 0.001
R6_4 193 192 0.001
R6_5 192 191 0.001
R6_6 191 194 0.001
R6_7 184 185 0.001
R6_8 194 196 0.2
C6_81 194 273 7.7e-16
C6_82 196 273 7.7e-16
R6_9 192 194 0.2
C6_91 192 273 7e-16
C6_92 194 273 7e-16
R6_10 185 192 1
C6_101 185 273 2.8e-15
C6_102 192 273 2.8e-15
R6_11 190 193 1.5
C6_111 190 273 7.2e-15
C6_112 193 273 7.2e-15
R6_12 189 195 0.5
C6_121 189 273 1.47e-15
C6_122 195 273 1.47e-15
R6_13 186 189 0.7
C6_131 186 273 2.1e-15
C6_132 189 273 2.1e-15
R6_14 183 187 500
C6_141 183 273 1.5e-15
C6_142 187 273 1.5e-15
R5_1 199 214 0.001
R5_2 200 223 0.001
R5_3 208 220 0.001
R5_4 200 209 0.001
R5_5 200 212 0.001
R5_6 200 201 0.001
R5_7 202 224 0.001
R5_8 203 228 0.001
R5_9 204 238 0.001
R5_10 210 232 0.001
R5_11 204 211 0.001
R5_12 204 213 0.001
R5_13 204 205 0.001
R5_14 206 240 0.001
R5_15 207 244 0.001
R5_16 243 247 0.001
C5_161 243 273 1.32e-15
C5_162 247 273 1.32e-15
R5_17 244 243 0.1
C5_171 244 273 1.44e-15
C5_172 243 273 1.44e-15
R5_18 245 244 0.001
C5_181 245 273 8.4e-16
C5_182 244 273 8.4e-16
R5_19 246 245 0.001
C5_191 246 273 2.4e-16
C5_192 245 273 2.4e-16
R5_20 239 246 0.001
C5_201 239 273 1.08e-15
C5_202 246 273 1.08e-15
R5_21 240 239 0.1
C5_211 240 273 1.44e-15
C5_212 239 273 1.44e-15
R5_22 241 240 0.001
C5_221 241 273 8.4e-16
C5_222 240 273 8.4e-16
R5_23 213 238 0.3
C5_231 213 273 9.8e-16
C5_232 238 273 9.8e-16
R5_24 211 213 0.2
C5_241 211 273 7e-16
C5_242 213 273 7e-16
R5_25 205 211 0.2
C5_251 205 273 7e-16
C5_252 211 273 7e-16
R5_26 242 241 0.001
C5_261 242 273 2.4e-16
C5_262 241 273 2.4e-16
R5_27 238 242 0.1
C5_271 238 273 2.28e-15
C5_272 242 273 2.28e-15
R5_28 235 238 0.1
C5_281 235 273 2.4e-15
C5_282 238 273 2.4e-15
R5_29 236 235 0.001
C5_291 236 273 1.2e-15
C5_292 235 273 1.2e-15
R5_30 237 236 0.001
C5_301 237 273 1.2e-15
C5_302 236 273 1.2e-15
R5_31 232 237 0.1
C5_311 232 273 1.44e-15
C5_312 237 273 1.44e-15
R5_32 233 232 0.1
C5_321 233 273 2.04e-15
C5_322 232 273 2.04e-15
R5_33 234 233 0.001
C5_331 234 273 2.4e-16
C5_332 233 273 2.4e-16
R5_34 231 234 0.001
C5_341 231 273 1.08e-15
C5_342 234 273 1.08e-15
R5_35 228 231 0.1
C5_351 228 273 1.44e-15
C5_352 231 273 1.44e-15
R5_36 229 228 0.001
C5_361 229 273 8.4e-16
C5_362 228 273 8.4e-16
R5_37 230 229 0.001
C5_371 230 273 2.4e-16
C5_372 229 273 2.4e-16
R5_38 227 230 0.001
C5_381 227 273 1.08e-15
C5_382 230 273 1.08e-15
R5_39 224 227 0.1
C5_391 224 273 1.44e-15
C5_392 227 273 1.44e-15
R5_40 225 224 0.001
C5_401 225 273 8.4e-16
C5_402 224 273 8.4e-16
R5_41 212 223 0.3
C5_411 212 273 9.8e-16
C5_412 223 273 9.8e-16
R5_42 209 212 0.2
C5_421 209 273 7e-16
C5_422 212 273 7e-16
R5_43 201 209 0.2
C5_431 201 273 7e-16
C5_432 209 273 7e-16
R5_44 226 225 0.001
C5_441 226 273 2.4e-16
C5_442 225 273 2.4e-16
R5_45 223 226 0.1
C5_451 223 273 2.28e-15
C5_452 226 273 2.28e-15
R5_46 221 223 0.1
C5_461 221 273 2.4e-15
C5_462 223 273 2.4e-15
R5_47 222 221 0.001
C5_471 222 273 1.2e-15
C5_472 221 273 1.2e-15
R5_48 219 222 0.001
C5_481 219 273 1.2e-15
C5_482 222 273 1.2e-15
R5_49 220 219 0.1
C5_491 220 273 1.44e-15
C5_492 219 273 1.44e-15
R5_50 216 220 0.1
C5_501 216 273 2.04e-15
C5_502 220 273 2.04e-15
R5_51 217 216 0.001
C5_511 217 273 2.4e-16
C5_512 216 273 2.4e-16
R5_52 215 217 0.001
C5_521 215 273 1.08e-15
C5_522 217 273 1.08e-15
R5_53 214 215 0.1
C5_531 214 273 1.5e-15
C5_532 215 273 1.5e-15
R5_54 218 214 0.001
C5_541 218 273 1.02e-15
C5_542 214 273 1.02e-15
R3_1 253 254 0.001
R3_2 262 263 0.001
R3_3 268 267 0.001
R3_4 262 264 0.001
R3_5 270 269 0.001
R3_6 260 259 0.001
R3_7 258 265 850
C3_71 258 273 2.625e-15
C3_72 265 273 2.625e-15
R3_8 255 258 750
C3_81 255 273 2.25e-15
C3_82 258 273 2.25e-15
R3_9 256 261 750
C3_91 256 273 2.25e-15
C3_92 261 273 2.25e-15
R3_10 259 266 850
C3_101 259 273 2.625e-15
C3_102 266 273 2.625e-15
R3_11 259 261 450
C3_111 259 273 1.35e-15
C3_112 261 273 1.35e-15
R3_12 258 259 450
C3_121 258 273 1.35e-15
C3_122 259 273 1.35e-15
R3_13 260 269 1
C3_131 260 273 2.8e-15
C3_132 269 273 2.8e-15
R3_14 257 260 0.2
C3_141 257 273 7.7e-16
C3_142 260 273 7.7e-16
R3_15 268 270 0.5
C3_151 268 273 2.4e-15
C3_152 270 273 2.4e-15
R3_16 263 267 0.2
C3_161 263 273 7e-16
C3_162 267 273 7e-16
R3_17 264 263 0.2
C3_171 264 273 7e-16
C3_172 263 273 7e-16
R3_18 254 264 1
C3_181 254 273 2.8e-15
C3_182 264 273 2.8e-15
R2_1 296 277 0.001
R2_2 297 278 0.001
R2_3 301 281 0.001
R2_4 297 305 0.001
R2_5 300 273 0.001
R2_6 302 282 0.001
R2_7 299 288 0.001
R2_8 298 285 0.001
R2_9 303 289 0.001
R2_10 299 306 0.001
R2_11 304 292 0.001
R2_12 292 294 0.1
C2_121 292 273 2.76e-15
C2_122 294 273 2.76e-15
R2_13 293 292 0.001
C2_131 293 273 8.4e-16
C2_132 292 273 8.4e-16
R2_14 288 306 0.3
C2_141 288 273 9.8e-16
C2_142 306 273 9.8e-16
R2_15 295 293 0.001
C2_151 295 273 2.4e-16
C2_152 293 273 2.4e-16
R2_16 289 295 0.1
C2_161 289 273 2.52e-15
C2_162 295 273 2.52e-15
R2_17 290 289 0.001
C2_171 290 273 8.4e-16
C2_172 289 273 8.4e-16
R2_18 291 290 0.001
C2_181 291 273 2.4e-16
C2_182 290 273 2.4e-16
R2_19 288 291 0.1
C2_191 288 273 2.28e-15
C2_192 291 273 2.28e-15
R2_20 285 288 0.4
C2_201 285 273 6.24e-15
C2_202 288 273 6.24e-15
R2_21 286 285 0.1
C2_211 286 273 2.04e-15
C2_212 285 273 2.04e-15
R2_22 287 286 0.001
C2_221 287 273 2.4e-16
C2_222 286 273 2.4e-16
R2_23 282 287 0.1
C2_231 282 273 2.52e-15
C2_232 287 273 2.52e-15
R2_24 283 282 0.001
C2_241 283 273 8.4e-16
C2_242 282 273 8.4e-16
R2_25 273 274 0.1
C2_251 273 273 2.58e-15
C2_252 274 273 2.58e-15
R2_26 276 273 0.001
C2_261 276 273 1.02e-15
C2_262 273 273 1.02e-15
R2_27 278 305 0.3
C2_271 278 273 9.8e-16
C2_272 305 273 9.8e-16
R2_28 284 283 0.001
C2_281 284 273 2.4e-16
C2_282 283 273 2.4e-16
R2_29 281 284 0.1
C2_291 281 273 2.52e-15
C2_292 284 273 2.52e-15
R2_30 279 281 0.001
C2_301 279 273 8.4e-16
C2_302 281 273 8.4e-16
R2_31 280 279 0.001
C2_311 280 273 2.4e-16
C2_312 279 273 2.4e-16
R2_32 278 280 0.1
C2_321 278 273 2.28e-15
C2_322 280 273 2.28e-15
R2_33 277 278 0.4
C2_331 277 273 6.24e-15
C2_332 278 273 6.24e-15
R2_34 275 277 0.1
C2_341 275 273 2.04e-15
C2_342 277 273 2.04e-15
R2_35 274 275 0.001
C2_351 274 273 2.4e-16
C2_352 275 273 2.4e-16
R1_1 309 310 0.001
R1_2 311 312 0.001
R1_3 316 319 0.001
R1_4 316 317 0.001
R1_5 315 314 0.001
R1_6 315 318 500
C1_61 315 273 1.575e-15
C1_62 318 273 1.575e-15
R1_7 313 314 1.7
C1_71 313 273 1.955e-15
C1_72 314 273 1.955e-15
R1_8 317 319 0.5
C1_81 317 273 5.75e-16
C1_82 319 273 5.75e-16
R1_9 310 317 2.5
C1_91 310 273 2.875e-15
C1_92 317 273 2.875e-15
R1_10 312 313 0.9
C1_101 312 273 1.035e-15
C1_102 313 273 1.035e-15
R1_11 310 312 1.3
C1_111 310 273 1.495e-15
C1_112 312 273 1.495e-15
.ends flipflop

