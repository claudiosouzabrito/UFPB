.include biel7.spi

V1 20 30 1.8V
V2 10 30 pulse (0V 1.8V 10ns 1ps 1ps 10ns 20ns)
V3 30 0 DC 0

x1 10 20 30 40 biel7
x2 40 20 30 42 biel7
x3 40 20 30 44 biel7
x4 40 20 30 46 biel7
x5 40 20 30 48 biel7

.model tp pmos level = 54
.model tn nmos level = 54

.tran 0.001ns 30ns
.end
