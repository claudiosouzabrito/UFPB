* Spice description of flipflopphi
* Spice driver version 224949768
* Date ( dd/mm/yyyy hh:mm:ss ): 20/08/2019 at 15:14:34

* INTERF d ph0 ph1 q vdd vss 


.subckt flipflopphi 218 230 58 43 149 254 
* NET 13 = latch2.inv1.nq
* NET 43 = q
* NET 58 = ph1
* NET 61 = latch2.mux.i0
* NET 149 = vdd
* NET 152 = latch1.mux.q
* NET 179 = latch1.inv1.nq
* NET 196 = latch1.mux.i0
* NET 218 = d
* NET 230 = ph0
* NET 254 = vss
Mtr_00032 109 85 39 149 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00031 1 169 109 149 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00030 99 56 115 149 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00029 4 57 87 149 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00028 87 101 1 149 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00027 115 66 4 149 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00026 20 41 111 149 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00025 69 19 112 149 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00024 105 290 167 149 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00023 10 216 105 149 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00022 246 228 113 149 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00021 7 229 292 149 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00020 292 248 10 149 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00019 113 201 7 149 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00018 186 166 107 149 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00017 204 185 108 149 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00016 278 154 30 254 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00015 30 51 80 254 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00014 277 49 92 254 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00013 80 94 77 254 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00012 77 61 277 254 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00011 33 81 278 254 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00010 279 36 13 254 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00009 280 16 62 254 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00008 274 212 236 254 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00007 236 223 285 254 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00006 273 221 239 254 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00005 285 241 233 254 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00004 233 196 273 254 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00003 152 286 274 254 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00002 275 153 179 254 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00001 276 182 197 254 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
R19_1 13 14 0.001
R19_2 20 22 0.001
R19_3 23 22 0.001
R19_4 20 21 0.001
R19_5 25 24 0.001
R19_6 18 17 0.001
R19_7 18 19 600
C19_71 18 254 1.875e-15
C19_72 19 254 1.875e-15
R19_8 16 18 500
C19_81 16 254 1.5e-15
C19_82 18 254 1.5e-15
R19_9 24 27 0.2
C19_91 24 254 7.7e-16
C19_92 27 254 7.7e-16
R19_10 17 24 0.7
C19_101 17 254 2.1e-15
C19_102 24 254 2.1e-15
R19_11 15 17 0.5
C19_111 15 254 1.47e-15
C19_112 17 254 1.47e-15
R19_12 23 25 0.25
C19_121 23 254 1.2e-15
C19_122 25 254 1.2e-15
R19_13 22 26 0.2
C19_131 22 254 7.7e-16
C19_132 26 254 7.7e-16
R19_14 21 22 0.2
C19_141 21 254 7e-16
C19_142 22 254 7e-16
R19_15 14 21 1
C19_151 14 254 2.8e-15
C19_152 21 254 2.8e-15
R17_1 33 34 0.001
R17_2 39 42 0.001
R17_3 39 43 0.001
R17_4 44 43 0.001
R17_5 39 40 0.001
R17_6 46 45 0.001
R17_7 38 37 0.001
R17_8 38 41 600
C17_81 38 254 1.875e-15
C17_82 41 254 1.875e-15
R17_9 36 38 500
C17_91 36 254 1.5e-15
C17_92 38 254 1.5e-15
R17_10 37 45 1
C17_101 37 254 2.8e-15
C17_102 45 254 2.8e-15
R17_11 35 37 0.5
C17_111 35 254 1.47e-15
C17_112 37 254 1.47e-15
R17_12 44 46 0.25
C17_121 44 254 1.2e-15
C17_122 46 254 1.2e-15
R17_13 42 43 0.2
C17_131 42 254 7e-16
C17_132 43 254 7e-16
R17_14 40 42 0.2
C17_141 40 254 7e-16
C17_142 42 254 7e-16
R17_15 34 40 1
C17_151 34 254 2.8e-15
C17_152 40 254 2.8e-15
R16_1 54 53 0.001
R16_2 53 58 1
C16_21 53 254 2.8e-15
C16_22 58 254 2.8e-15
R16_3 50 53 0.2
C16_31 50 254 7.7e-16
C16_32 53 254 7.7e-16
R16_4 54 57 850
C16_41 54 254 2.625e-15
C16_42 57 254 2.625e-15
R16_5 51 55 750
C16_51 51 254 2.25e-15
C16_52 55 254 2.25e-15
R16_6 54 55 450
C16_61 54 254 1.35e-15
C16_62 55 254 1.35e-15
R16_7 52 54 450
C16_71 52 254 1.35e-15
C16_72 54 254 1.35e-15
R16_8 52 56 850
C16_81 52 254 2.625e-15
C16_82 56 254 2.625e-15
R16_9 49 52 750
C16_91 49 254 2.25e-15
C16_92 52 254 2.25e-15
R15_1 65 64 0.001
R15_2 66 67 0.001
R15_3 68 67 0.001
R15_4 71 70 0.001
R15_5 70 69 0.001
R15_6 69 72 0.001
R15_7 62 63 0.001
R15_8 72 74 0.2
C15_81 72 254 7.7e-16
C15_82 74 254 7.7e-16
R15_9 70 72 0.2
C15_91 70 254 7e-16
C15_92 72 254 7e-16
R15_10 63 70 1
C15_101 63 254 2.8e-15
C15_102 70 254 2.8e-15
R15_11 68 71 1.5
C15_111 68 254 7.2e-15
C15_112 71 254 7.2e-15
R15_12 67 73 0.5
C15_121 67 254 1.47e-15
C15_122 73 254 1.47e-15
R15_13 64 67 0.7
C15_131 64 254 2.1e-15
C15_132 67 254 2.1e-15
R15_14 61 65 500
C15_141 61 254 1.5e-15
C15_142 65 254 1.5e-15
R13_1 80 82 0.001
R13_2 87 88 0.001
R13_3 87 89 0.001
R13_4 84 83 0.001
R13_5 86 85 700
C13_51 86 254 2.175e-15
C13_52 85 254 2.175e-15
R13_6 81 86 750
C13_61 81 254 2.325e-15
C13_62 86 254 2.325e-15
R13_7 84 86 900
C13_71 84 254 2.7e-15
C13_72 86 254 2.7e-15
R13_8 88 89 0.5
C13_81 88 254 5.75e-16
C13_82 89 254 5.75e-16
R13_9 83 88 1.1
C13_91 83 254 1.265e-15
C13_92 88 254 1.265e-15
R13_10 82 83 0.9
C13_101 82 254 1.035e-15
C13_102 83 254 1.035e-15
R12_1 92 93 0.001
R12_2 99 102 0.001
R12_3 99 100 0.001
R12_4 94 95 0.001
R12_5 98 97 0.001
R12_6 98 101 500
C12_61 98 254 1.575e-15
C12_62 101 254 1.575e-15
R12_7 96 97 1.7
C12_71 96 254 1.955e-15
C12_72 97 254 1.955e-15
R12_8 95 96 0.9
C12_81 95 254 1.035e-15
C12_82 96 254 1.035e-15
R12_9 93 95 1.3
C12_91 93 254 1.495e-15
C12_92 95 254 1.495e-15
R12_10 100 102 0.5
C12_101 100 254 5.75e-16
C12_102 102 254 5.75e-16
R12_11 93 100 2.5
C12_111 93 254 2.875e-15
C12_112 100 254 2.875e-15
R11_1 105 114 0.001
R11_2 105 117 0.001
R11_3 105 124 0.001
R11_4 105 106 0.001
R11_5 113 119 0.001
R11_6 107 127 0.001
R11_7 108 131 0.001
R11_8 109 139 0.001
R11_9 115 134 0.001
R11_10 109 116 0.001
R11_11 109 118 0.001
R11_12 109 110 0.001
R11_13 111 142 0.001
R11_14 112 146 0.001
R11_15 145 148 0.001
C11_151 145 254 1.32e-15
C11_152 148 254 1.32e-15
R11_16 146 145 0.1
C11_161 146 254 1.44e-15
C11_162 145 254 1.44e-15
R11_17 147 146 0.001
C11_171 147 254 8.4e-16
C11_172 146 254 8.4e-16
R11_18 143 147 0.001
C11_181 143 254 2.4e-16
C11_182 147 254 2.4e-16
R11_19 141 143 0.001
C11_191 141 254 1.08e-15
C11_192 143 254 1.08e-15
R11_20 142 141 0.1
C11_201 142 254 1.44e-15
C11_202 141 254 1.44e-15
R11_21 144 142 0.001
C11_211 144 254 8.4e-16
C11_212 142 254 8.4e-16
R11_22 118 139 0.3
C11_221 118 254 9.8e-16
C11_222 139 254 9.8e-16
R11_23 116 118 0.2
C11_231 116 254 7e-16
C11_232 118 254 7e-16
R11_24 110 116 0.2
C11_241 110 254 7e-16
C11_242 116 254 7e-16
R11_25 140 144 0.001
C11_251 140 254 2.4e-16
C11_252 144 254 2.4e-16
R11_26 139 140 0.1
C11_261 139 254 2.28e-15
C11_262 140 254 2.28e-15
R11_27 137 139 0.1
C11_271 137 254 2.4e-15
C11_272 139 254 2.4e-15
R11_28 138 137 0.001
C11_281 138 254 1.2e-15
C11_282 137 254 1.2e-15
R11_29 135 138 0.001
C11_291 135 254 1.2e-15
C11_292 138 254 1.2e-15
R11_30 134 135 0.1
C11_301 134 254 1.44e-15
C11_302 135 254 1.44e-15
R11_31 136 134 0.1
C11_311 136 254 2.04e-15
C11_312 134 254 2.04e-15
R11_32 132 136 0.001
C11_321 132 254 2.4e-16
C11_322 136 254 2.4e-16
R11_33 130 132 0.001
C11_331 130 254 1.08e-15
C11_332 132 254 1.08e-15
R11_34 131 130 0.1
C11_341 131 254 1.44e-15
C11_342 130 254 1.44e-15
R11_35 133 131 0.001
C11_351 133 254 8.4e-16
C11_352 131 254 8.4e-16
R11_36 128 133 0.001
C11_361 128 254 2.4e-16
C11_362 133 254 2.4e-16
R11_37 126 128 0.001
C11_371 126 254 1.08e-15
C11_372 128 254 1.08e-15
R11_38 127 126 0.1
C11_381 127 254 1.44e-15
C11_382 126 254 1.44e-15
R11_39 129 127 0.001
C11_391 129 254 8.4e-16
C11_392 127 254 8.4e-16
R11_40 125 129 0.001
C11_401 125 254 2.4e-16
C11_402 129 254 2.4e-16
R11_41 124 125 0.1
C11_411 124 254 2.28e-15
C11_412 125 254 2.28e-15
R11_42 124 149 0.001
C11_421 124 254 4.8e-16
C11_422 149 254 4.8e-16
R11_43 123 149 0.1
C11_431 123 254 1.92e-15
C11_432 149 254 1.92e-15
R11_44 122 123 0.001
C11_441 122 254 1.2e-15
C11_442 123 254 1.2e-15
R11_45 120 122 0.001
C11_451 120 254 1.2e-15
C11_452 122 254 1.2e-15
R11_46 119 120 0.1
C11_461 119 254 1.44e-15
C11_462 120 254 1.44e-15
R11_47 121 119 0.1
C11_471 121 254 2.28e-15
C11_472 119 254 2.28e-15
R11_48 117 124 0.3
C11_481 117 254 9.8e-16
C11_482 124 254 9.8e-16
R11_49 114 117 0.2
C11_491 114 254 7e-16
C11_492 117 254 7e-16
R11_50 106 114 0.2
C11_501 106 254 7e-16
C11_502 114 254 7e-16
R10_1 152 155 0.001
R10_2 167 171 0.001
R10_3 167 172 0.001
R10_4 173 172 0.001
R10_5 167 168 0.001
R10_6 161 160 0.001
R10_7 175 174 0.001
R10_8 165 164 0.001
R10_9 163 162 0.001
R10_10 158 157 0.001
R10_11 169 170 0.001
R10_12 154 158 500
C10_121 154 254 1.5e-15
C10_122 158 254 1.5e-15
R10_13 163 166 600
C10_131 163 254 1.875e-15
C10_132 166 254 1.875e-15
R10_14 153 163 500
C10_141 153 254 1.5e-15
C10_142 163 254 1.5e-15
R10_15 170 176 0.5
C10_151 170 254 1.47e-15
C10_152 176 254 1.47e-15
R10_16 164 170 0.5
C10_161 164 254 1.4e-15
C10_162 170 254 1.4e-15
R10_17 157 164 0.2
C10_171 157 254 7e-16
C10_172 164 254 7e-16
R10_18 159 157 0.2
C10_181 159 254 7.7e-16
C10_182 157 254 7.7e-16
R10_19 162 174 1
C10_191 162 254 2.8e-15
C10_192 174 254 2.8e-15
R10_20 156 162 0.5
C10_201 156 254 1.47e-15
C10_202 162 254 1.47e-15
R10_21 161 165 1.6
C10_211 161 254 7.8e-15
C10_212 165 254 7.8e-15
R10_22 173 175 0.25
C10_221 173 254 1.2e-15
C10_222 175 254 1.2e-15
R10_23 171 172 0.2
C10_231 171 254 7e-16
C10_232 172 254 7e-16
R10_24 168 171 0.2
C10_241 168 254 7e-16
C10_242 171 254 7e-16
R10_25 160 168 0.5
C10_251 160 254 1.4e-15
C10_252 168 254 1.4e-15
R10_26 155 160 0.5
C10_261 155 254 1.4e-15
C10_262 160 254 1.4e-15
R9_1 179 180 0.001
R9_2 186 188 0.001
R9_3 189 188 0.001
R9_4 186 187 0.001
R9_5 191 190 0.001
R9_6 184 183 0.001
R9_7 184 185 600
C9_71 184 254 1.875e-15
C9_72 185 254 1.875e-15
R9_8 182 184 500
C9_81 182 254 1.5e-15
C9_82 184 254 1.5e-15
R9_9 190 193 0.2
C9_91 190 254 7.7e-16
C9_92 193 254 7.7e-16
R9_10 183 190 0.7
C9_101 183 254 2.1e-15
C9_102 190 254 2.1e-15
R9_11 181 183 0.5
C9_111 181 254 1.47e-15
C9_112 183 254 1.47e-15
R9_12 189 191 0.25
C9_121 189 254 1.2e-15
C9_122 191 254 1.2e-15
R9_13 188 192 0.2
C9_131 188 254 7.7e-16
C9_132 192 254 7.7e-16
R9_14 187 188 0.2
C9_141 187 254 7e-16
C9_142 188 254 7e-16
R9_15 180 187 1
C9_151 180 254 2.8e-15
C9_152 187 254 2.8e-15
R8_1 200 199 0.001
R8_2 201 202 0.001
R8_3 203 202 0.001
R8_4 206 205 0.001
R8_5 205 204 0.001
R8_6 204 207 0.001
R8_7 197 198 0.001
R8_8 207 209 0.2
C8_81 207 254 7.7e-16
C8_82 209 254 7.7e-16
R8_9 205 207 0.2
C8_91 205 254 7e-16
C8_92 207 254 7e-16
R8_10 198 205 1
C8_101 198 254 2.8e-15
C8_102 205 254 2.8e-15
R8_11 203 206 1.5
C8_111 203 254 7.2e-15
C8_112 206 254 7.2e-15
R8_12 202 208 0.5
C8_121 202 254 1.47e-15
C8_122 208 254 1.47e-15
R8_13 199 202 0.7
C8_131 199 254 2.1e-15
C8_132 202 254 2.1e-15
R8_14 196 200 500
C8_141 196 254 1.5e-15
C8_142 200 254 1.5e-15
R7_1 213 214 0.001
R7_2 216 217 0.001
R7_3 217 218 0.5
C7_31 217 254 1.4e-15
C7_32 218 254 1.4e-15
R7_4 214 217 0.7
C7_41 214 254 2.1e-15
C7_42 217 254 2.1e-15
R7_5 215 214 0.2
C7_51 215 254 7.7e-16
C7_52 214 254 7.7e-16
R7_6 212 213 500
C7_61 212 254 1.5e-15
C7_62 213 254 1.5e-15
R6_1 226 225 0.001
R6_2 225 230 1
C6_21 225 254 2.8e-15
C6_22 230 254 2.8e-15
R6_3 222 225 0.2
C6_31 222 254 7.7e-16
C6_32 225 254 7.7e-16
R6_4 226 229 850
C6_41 226 254 2.625e-15
C6_42 229 254 2.625e-15
R6_5 224 228 850
C6_51 224 254 2.625e-15
C6_52 228 254 2.625e-15
R6_6 221 224 750
C6_61 221 254 2.25e-15
C6_62 224 254 2.25e-15
R6_7 226 227 450
C6_71 226 254 1.35e-15
C6_72 227 254 1.35e-15
R6_8 224 226 450
C6_81 224 254 1.35e-15
C6_82 226 254 1.35e-15
R6_9 223 227 750
C6_91 223 254 2.25e-15
C6_92 227 254 2.25e-15
R3_1 239 240 0.001
R3_2 246 249 0.001
R3_3 246 247 0.001
R3_4 241 242 0.001
R3_5 245 244 0.001
R3_6 245 248 500
C3_61 245 254 1.575e-15
C3_62 248 254 1.575e-15
R3_7 243 244 1.7
C3_71 243 254 1.955e-15
C3_72 244 254 1.955e-15
R3_8 242 243 0.9
C3_81 242 254 1.035e-15
C3_82 243 254 1.035e-15
R3_9 240 242 1.3
C3_91 240 254 1.495e-15
C3_92 242 254 1.495e-15
R3_10 247 249 0.5
C3_101 247 254 5.75e-16
C3_102 249 254 5.75e-16
R3_11 240 247 2.5
C3_111 240 254 2.875e-15
C3_112 247 254 2.875e-15
R2_1 273 252 0.001
R2_2 274 255 0.001
R2_3 275 256 0.001
R2_4 274 281 0.001
R2_5 276 257 0.001
R2_6 278 265 0.001
R2_7 277 262 0.001
R2_8 278 282 0.001
R2_9 279 266 0.001
R2_10 280 269 0.001
R2_11 269 272 0.1
C2_111 269 254 2.76e-15
C2_112 272 254 2.76e-15
R2_12 270 269 0.001
C2_121 270 254 8.4e-16
C2_122 269 254 8.4e-16
R2_13 271 270 0.001
C2_131 271 254 2.4e-16
C2_132 270 254 2.4e-16
R2_14 266 271 0.1
C2_141 266 254 2.52e-15
C2_142 271 254 2.52e-15
R2_15 267 266 0.001
C2_151 267 254 8.4e-16
C2_152 266 254 8.4e-16
R2_16 265 282 0.3
C2_161 265 254 9.8e-16
C2_162 282 254 9.8e-16
R2_17 268 267 0.001
C2_171 268 254 2.4e-16
C2_172 267 254 2.4e-16
R2_18 265 268 0.1
C2_181 265 254 2.28e-15
C2_182 268 254 2.28e-15
R2_19 262 265 0.4
C2_191 262 254 6.24e-15
C2_192 265 254 6.24e-15
R2_20 263 262 0.1
C2_201 263 254 2.04e-15
C2_202 262 254 2.04e-15
R2_21 264 263 0.001
C2_211 264 254 2.4e-16
C2_212 263 254 2.4e-16
R2_22 257 264 0.1
C2_221 257 254 2.52e-15
C2_222 264 254 2.52e-15
R2_23 258 257 0.001
C2_231 258 254 8.4e-16
C2_232 257 254 8.4e-16
R2_24 255 281 0.3
C2_241 255 254 9.8e-16
C2_242 281 254 9.8e-16
R2_25 259 258 0.001
C2_251 259 254 2.4e-16
C2_252 258 254 2.4e-16
R2_26 256 259 0.1
C2_261 256 254 2.52e-15
C2_262 259 254 2.52e-15
R2_27 260 256 0.001
C2_271 260 254 8.4e-16
C2_272 256 254 8.4e-16
R2_28 261 260 0.001
C2_281 261 254 2.4e-16
C2_282 260 254 2.4e-16
R2_29 254 261 0.1
C2_291 254 254 1.8e-15
C2_292 261 254 1.8e-15
R2_30 255 254 0.001
C2_301 255 254 4.8e-16
C2_302 254 254 4.8e-16
R2_31 252 255 0.4
C2_311 252 254 6.24e-15
C2_312 255 254 6.24e-15
R2_32 253 252 0.1
C2_321 253 254 2.28e-15
C2_322 252 254 2.28e-15
R1_1 285 287 0.001
R1_2 292 293 0.001
R1_3 292 294 0.001
R1_4 289 288 0.001
R1_5 291 290 700
C1_51 291 254 2.175e-15
C1_52 290 254 2.175e-15
R1_6 286 291 750
C1_61 286 254 2.325e-15
C1_62 291 254 2.325e-15
R1_7 289 291 900
C1_71 289 254 2.7e-15
C1_72 291 254 2.7e-15
R1_8 293 294 0.5
C1_81 293 254 5.75e-16
C1_82 294 254 5.75e-16
R1_9 288 293 1.1
C1_91 288 254 1.265e-15
C1_92 293 254 1.265e-15
R1_10 287 288 0.9
C1_101 287 254 1.035e-15
C1_102 288 254 1.035e-15
.ends flipflopphi

