* Spice description of gordo
* Spice driver version -360483320
* Date ( dd/mm/yyyy hh:mm:ss ):  9/07/2019 at 16:07:13

* INTERF a vdd vss y 


.subckt gordo 3 13 21 30 
* NET 3 = a
* NET 13 = vdd
* NET 21 = vss
* NET 30 = y
Mtr_00002 10 5 29 13 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_00001 18 2 26 21 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
R4_1 4 3 0.001
R4_2 6 5 650
C4_21 6 21 1.95e-15
C4_22 5 21 1.95e-15
R4_3 2 6 450
C4_31 2 21 1.425e-15
C4_32 6 21 1.425e-15
R4_4 3 7 0.9
C4_41 3 21 2.73e-15
C4_42 7 21 2.73e-15
R4_5 1 3 0.4
C4_51 1 21 1.33e-15
C4_52 3 21 1.33e-15
R4_6 4 6 200
C4_61 4 21 6e-16
C4_62 6 21 6e-16
R3_1 10 11 0.001
R3_2 14 15 0.001
C3_21 14 21 6e-16
C3_22 15 21 6e-16
R3_3 14 13 0.001
C3_31 14 21 1.2e-15
C3_32 13 21 1.2e-15
R3_4 11 13 0.001
C3_41 11 21 1.2e-15
C3_42 13 21 1.2e-15
R3_5 12 11 0.001
C3_51 12 21 8.4e-16
C3_52 11 21 8.4e-16
R2_1 18 19 0.001
R2_2 22 23 0.001
C2_21 22 21 6e-16
C2_22 23 21 6e-16
R2_3 22 21 0.001
C2_31 22 21 1.2e-15
C2_32 21 21 1.2e-15
R2_4 19 21 0.001
C2_41 19 21 1.2e-15
C2_42 21 21 1.2e-15
R2_5 20 19 0.001
C2_51 20 21 8.4e-16
C2_52 19 21 8.4e-16
R1_1 26 27 0.001
R1_2 29 31 0.001
R1_3 31 32 0.1
C1_31 31 21 4.9e-16
C1_32 32 21 4.9e-16
R1_4 30 31 0.8
C1_41 30 21 2.24e-15
C1_42 31 21 2.24e-15
R1_5 27 30 0.3
C1_51 27 21 9.8e-16
C1_52 30 21 9.8e-16
R1_6 28 27 0.1
C1_61 28 21 3.5e-16
C1_62 27 21 3.5e-16
.ends gordo

