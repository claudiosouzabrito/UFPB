* Spice description of gordo2
* Spice driver version -796658168
* Date ( dd/mm/yyyy hh:mm:ss ): 11/07/2019 at  0:28:43

* INTERF a vdd vss y 


.subckt gordo2 4 15 32 24 
* NET 4 = a
* NET 15 = vdd
* NET 24 = y
* NET 32 = vss
Mtr_00002 12 6 23 15 tp L=1U W=19U AS=38P AD=38P PS=42U PD=42U 
Mtr_00001 29 2 20 32 tn L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
R4_1 5 4 0.001
R4_2 2 3 300
C4_21 2 32 9e-16
C4_22 3 32 9e-16
R4_3 8 6 650
C4_31 8 32 1.95e-15
C4_32 6 32 1.95e-15
R4_4 7 8 50
C4_41 7 32 2.25e-16
C4_42 8 32 2.25e-16
R4_5 3 7 150
C4_51 3 32 4.5e-16
C4_52 7 32 4.5e-16
R4_6 4 9 0.9
C4_61 4 32 2.73e-15
C4_62 9 32 2.73e-15
R4_7 1 4 0.4
C4_71 1 32 1.33e-15
C4_72 4 32 1.33e-15
R4_8 5 8 200
C4_81 5 32 6e-16
C4_82 8 32 6e-16
R3_1 12 13 0.001
R3_2 16 17 0.001
C3_21 16 32 6e-16
C3_22 17 32 6e-16
R3_3 16 15 0.001
C3_31 16 32 1.2e-15
C3_32 15 32 1.2e-15
R3_4 13 15 0.001
C3_41 13 32 1.2e-15
C3_42 15 32 1.2e-15
R3_5 14 13 0.001
C3_51 14 32 8.4e-16
C3_52 13 32 8.4e-16
R2_1 20 21 0.001
R2_2 23 25 0.001
R2_3 25 26 0.1
C2_31 25 32 4.9e-16
C2_32 26 32 4.9e-16
R2_4 24 25 0.8
C2_41 24 32 2.24e-15
C2_42 25 32 2.24e-15
R2_5 21 24 0.4
C2_51 21 32 1.12e-15
C2_52 24 32 1.12e-15
R2_6 22 21 0.001
C2_61 22 32 2.1e-16
C2_62 21 32 2.1e-16
R1_1 29 30 0.001
R1_2 33 34 0.001
C1_21 33 32 6e-16
C1_22 34 32 6e-16
R1_3 33 32 0.001
C1_31 33 32 1.2e-15
C1_32 32 32 1.2e-15
R1_4 30 32 0.001
C1_41 30 32 1.2e-15
C1_42 32 32 1.2e-15
R1_5 31 30 0.001
C1_51 31 32 8.4e-16
C1_52 30 32 8.4e-16
.ends gordo2

