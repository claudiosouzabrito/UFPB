.include 2faseclk.spi

* INTERF clk q qb vdd vss vss
x1 10 40 41 20 30 30 2faseclk

v4 20 30 1.8V
v5 30 0 0V DC


v3 10 30 pulse(0 1.8 0ns 1ps 1ps 49ns 100ns)

.tran 0.01ns 400ns

.model tp pmos level=54
.model tn nmos level=54

.end 
