.include inversor5.spi

V1 20 30 1.8V
V2 10 30 pulse (0V 1.8V 10ns 1ps 1ps 10ns 20ns)
V3 30 0 DC 0

x1 10 20 30 40 inversor5
x2 40 20 30 41 inversor5
x3 40 20 30 42 inversor5
x4 40 20 30 43 inversor5
x5 40 20 30 44 inversor5

.model tp pmos level = 54
.model tn nmos level = 54

.tran 0.001ns 30ns
.end
