.include 2faseclk.spi
.include inv_x1.spi
.include flipflopphi.spi

* INTERF clk q qb vdd vss vss
x1        10 40 41 20 30 30 2faseclk

*INTERF i nq vdd vss
x2     40 42 20 30 inv_x1
x3     41 43 20 30 inv_x1 

* INTERF d ph0 ph1 q vdd vss 
x4       11 43 42 44 20 30 flipflopphi

v4 20 30 1.8V
v5 30 0 0V DC


v3 10 30 pulse(0 1.8 0ns 1ps 1ps 40ns 80ns)
v6 11 30 pulse(0 1.8 0ns 1ps 1ps 25ns 50ns)

.tran 0.01ns 400ns

.model tp pmos level=54
.model tn nmos level=54

.end 
