* Spice description of tiristorinversor
* Spice driver version -2022803960
* Date ( dd/mm/yyyy hh:mm:ss ): 30/07/2019 at 15:21:35

* INTERF a s vdd vss y 


.subckt tiristorinversor 13 31 45 77 6 
* NET 6 = y
* NET 13 = a
* NET 31 = s
* NET 45 = vdd
* NET 54 = inversor_1.nq
* NET 77 = vss
Mtr_00009 59 33 40 45 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00008 40 33 59 45 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00007 37 61 5 45 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00006 41 18 37 45 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00005 72 21 54 77 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00004 51 27 1 77 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00003 72 21 54 77 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00002 51 27 1 77 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00001 78 16 51 77 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
R8_1 1 2 0.001
R8_2 5 7 0.001
R8_3 7 9 0.2
C8_31 7 77 2.875e-16
C8_32 9 77 2.875e-16
R8_4 8 7 0.1
C8_41 8 77 1.725e-16
C8_42 7 77 1.725e-16
R8_5 10 8 0.1
C8_51 10 77 1.15e-16
C8_52 8 77 1.15e-16
R8_6 6 10 1
C8_61 6 77 1.2075e-15
C8_62 10 77 1.2075e-15
R8_7 3 6 0.9
C8_71 3 77 1.0925e-15
C8_72 6 77 1.0925e-15
R8_8 4 3 0.1
C8_81 4 77 1.15e-16
C8_82 3 77 1.15e-16
R8_9 2 4 0.1
C8_91 2 77 1.725e-16
C8_92 4 77 1.725e-16
R7_1 14 13 0.001
R7_2 13 17 1.5
C7_21 13 77 1.7825e-15
C7_22 17 77 1.7825e-15
R7_3 15 13 0.9
C7_31 15 77 1.0925e-15
C7_32 13 77 1.0925e-15
R7_4 14 18 550
C7_41 14 77 1.65e-15
C7_42 18 77 1.65e-15
R7_5 16 14 500
C7_51 16 77 1.5e-15
C7_52 14 77 1.5e-15
R6_1 32 31 0.001
R6_2 28 27 200
C6_21 28 77 6.75e-16
C6_22 27 77 6.75e-16
R6_3 29 28 50
C6_31 29 77 1.5e-16
C6_32 28 77 1.5e-16
R6_4 30 29 50
C6_41 30 77 2.25e-16
C6_42 29 77 2.25e-16
R6_5 25 30 700
C6_51 25 77 2.175e-15
C6_52 30 77 2.175e-15
R6_6 26 25 50
C6_61 26 77 1.5e-16
C6_62 25 77 1.5e-16
R6_7 23 26 300
C6_71 23 77 9.75e-16
C6_72 26 77 9.75e-16
R6_8 23 24 100
C6_81 23 77 3e-16
C6_82 24 77 3e-16
R6_9 31 34 1
C6_91 31 77 2.87e-15
C6_92 34 77 2.87e-15
R6_10 22 31 0.5
C6_101 22 77 1.47e-15
C6_102 31 77 1.47e-15
R6_11 21 24 400
C6_111 21 77 1.2e-15
C6_112 24 77 1.2e-15
R6_12 32 33 700
C6_121 32 77 2.1e-15
C6_122 33 77 2.1e-15
R6_13 21 32 450
C6_131 21 77 1.35e-15
C6_132 32 77 1.35e-15
R4_1 41 47 0.001
R4_2 40 42 0.001
R4_3 47 48 0.3
C4_31 47 77 4.92e-15
C4_32 48 77 4.92e-15
R4_4 45 47 0.1
C4_41 45 77 2.4e-15
C4_42 47 77 2.4e-15
R4_5 46 45 0.001
C4_51 46 77 1.2e-15
C4_52 45 77 1.2e-15
R4_6 42 46 0.1
C4_61 42 77 1.56e-15
C4_62 46 77 1.56e-15
R4_7 43 42 0.001
C4_71 43 77 9.6e-16
C4_72 42 77 9.6e-16
R4_8 44 43 0.001
C4_81 44 77 2.4e-16
C4_82 43 77 2.4e-16
R2_1 54 55 0.001
R2_2 59 62 0.001
R2_3 59 60 0.001
R2_4 57 56 0.001
R2_5 61 67 400
C2_51 61 77 1.275e-15
C2_52 67 77 1.275e-15
R2_6 68 69 50
C2_61 68 77 2.25e-16
C2_62 69 77 2.25e-16
R2_7 67 68 50
C2_71 67 77 1.5e-16
C2_72 68 77 1.5e-16
R2_8 65 69 700
C2_81 65 77 2.175e-15
C2_82 69 77 2.175e-15
R2_9 66 65 50
C2_91 66 77 1.5e-16
C2_92 65 77 1.5e-16
R2_10 64 66 300
C2_101 64 77 9.75e-16
C2_102 66 77 9.75e-16
R2_11 58 64 1200
C2_111 58 77 3.6e-15
C2_112 64 77 3.6e-15
R2_12 57 58 200
C2_121 57 77 6e-16
C2_122 58 77 6e-16
R2_13 62 63 0.2
C2_131 62 77 7.7e-16
C2_132 63 77 7.7e-16
R2_14 60 62 0.2
C2_141 60 77 7e-16
C2_142 62 77 7e-16
R2_15 56 60 0.5
C2_151 56 77 1.4e-15
C2_152 60 77 1.4e-15
R2_16 55 56 0.5
C2_161 55 77 1.4e-15
C2_162 56 77 1.4e-15
R1_1 72 73 0.001
R1_2 78 79 0.001
R1_3 79 80 0.3
C1_31 79 77 4.92e-15
C1_32 80 77 4.92e-15
R1_4 77 79 0.1
C1_41 77 77 2.4e-15
C1_42 79 77 2.4e-15
R1_5 76 75 0.001
C1_51 76 77 2.4e-16
C1_52 75 77 2.4e-16
R1_6 74 77 0.001
C1_61 74 77 1.2e-15
C1_62 77 77 1.2e-15
R1_7 73 74 0.1
C1_71 73 77 1.56e-15
C1_72 74 77 1.56e-15
R1_8 75 73 0.001
C1_81 75 77 9.6e-16
C1_82 73 77 9.6e-16
.ends tiristorinversor

