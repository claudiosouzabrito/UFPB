.include inv+fo4.spi
.include inversor5.spi
.include inv-gordo+fo4.spi
.include f04.spi

V1 20 30 1.8V
V2 10 30 pulse (0.0V 1.8V 10ns 1ps 1ps 10ns 20ns)
V3 30 0 DC 0

x2 10 20 30 40 inversor5
x1 10 20 30 41 inv+fo4
x3 10 20 30 42 inv-gordo+fo4
x4 10 20 30 43 inversor5
x5 10 20 30 43 inversor5
x6 43 20 30 f04

.model tp pmos level = 54
.model tn nmos level = 54

.tran 0.001ns 30ns
.end
