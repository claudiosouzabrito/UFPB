* Spice description of mux
* Spice driver version -63408632
* Date ( dd/mm/yyyy hh:mm:ss ):  1/08/2019 at 15:17:16

* INTERF d0 d1 s vdd-e vss-e y 


.subckt mux 18 11 81 107 113 35 
* NET 1 = tiristor2.inversor_1.vdd
* NET 11 = d1
* NET 18 = d0
* NET 35 = y
* NET 51 = tiristor2.inversor_1.vss
* NET 81 = s
* NET 107 = vdd-e
* NET 113 = vss-e
* NET 123 = tiristor1.inversor_1.nq
Mtr_00012 86 146 1 107 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00011 12 147 41 107 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00010 144 84 96 107 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00009 19 85 37 107 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00008 141 82 95 107 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00007 95 82 141 107 tp L=1U W=13U AS=26P AD=26P PS=30U PD=30U 
Mtr_00006 51 130 62 113 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00005 9 65 28 113 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00004 116 61 125 113 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00003 16 128 23 113 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00002 110 58 123 113 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00001 110 58 123 113 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
R9_1 1 2 0.001
R9_2 5 6 0.001
C9_21 5 113 6e-16
C9_22 6 113 6e-16
R9_3 4 5 0.001
C9_31 4 113 7.2e-16
C9_32 5 113 7.2e-16
R9_4 2 4 0.1
C9_41 2 113 1.44e-15
C9_42 4 113 1.44e-15
R9_5 3 2 0.001
C9_51 3 113 1.08e-15
C9_52 2 113 1.08e-15
R8_1 9 10 0.001
R8_2 12 13 0.001
R8_3 11 13 1.3
C8_31 11 113 1.495e-15
C8_32 13 113 1.495e-15
R8_4 10 11 1.2
C8_41 10 113 1.38e-15
C8_42 11 113 1.38e-15
R7_1 16 17 0.001
R7_2 19 20 0.001
R7_3 18 20 1.3
C7_31 18 113 1.495e-15
C7_32 20 113 1.495e-15
R7_4 17 18 1.2
C7_41 17 113 1.38e-15
C7_42 18 113 1.38e-15
R6_1 23 24 0.001
R6_2 34 33 0.001
R6_3 37 45 0.001
R6_4 36 35 0.001
R6_5 41 47 0.001
R6_6 28 29 0.001
R6_7 29 30 0.1
C6_71 29 113 1.725e-16
C6_72 30 113 1.725e-16
R6_8 32 29 0.2
C6_81 32 113 2.875e-16
C6_82 29 113 2.875e-16
R6_9 47 48 0.2
C6_91 47 113 2.875e-16
C6_92 48 113 2.875e-16
R6_10 42 47 0.1
C6_101 42 113 1.725e-16
C6_102 47 113 1.725e-16
R6_11 43 42 0.1
C6_111 43 113 1.15e-16
C6_112 42 113 1.15e-16
R6_12 35 43 1
C6_121 35 113 1.2075e-15
C6_122 43 113 1.2075e-15
R6_13 31 35 0.9
C6_131 31 113 1.0925e-15
C6_132 35 113 1.0925e-15
R6_14 30 31 0.1
C6_141 30 113 1.15e-16
C6_142 31 113 1.15e-16
R6_15 36 44 0.15
C6_151 36 113 8.4e-16
C6_152 44 113 8.4e-16
R6_16 38 44 0.75
C6_161 38 113 3.6e-15
C6_162 44 113 3.6e-15
R6_17 34 38 0.15
C6_171 34 113 8.4e-16
C6_172 38 113 8.4e-16
R6_18 45 46 0.2
C6_181 45 113 2.875e-16
C6_182 46 113 2.875e-16
R6_19 39 45 0.1
C6_191 39 113 1.725e-16
C6_192 45 113 1.725e-16
R6_20 40 39 0.1
C6_201 40 113 1.15e-16
C6_202 39 113 1.15e-16
R6_21 33 40 1
C6_211 33 113 1.2075e-15
C6_212 40 113 1.2075e-15
R6_22 25 33 0.9
C6_221 25 113 1.0925e-15
C6_222 33 113 1.0925e-15
R6_23 26 25 0.1
C6_231 26 113 1.15e-16
C6_232 25 113 1.15e-16
R6_24 24 26 0.1
C6_241 24 113 1.725e-16
C6_242 26 113 1.725e-16
R6_25 27 24 0.2
C6_251 27 113 2.875e-16
C6_252 24 113 2.875e-16
R5_1 51 52 0.001
R5_2 54 55 0.001
C5_21 54 113 6e-16
C5_22 55 113 6e-16
R5_3 52 54 0.1
C5_31 52 113 2.16e-15
C5_32 54 113 2.16e-15
R5_4 53 52 0.001
C5_41 53 113 1.08e-15
C5_42 52 113 1.08e-15
R4_1 73 72 0.001
R4_2 72 74 0.001
R4_3 83 81 0.001
R4_4 77 76 0.001
R4_5 76 78 0.001
R4_6 70 69 0.001
R4_7 86 88 0.001
R4_8 86 87 0.001
R4_9 62 63 0.001
R4_10 66 65 250
C4_101 66 113 7.5e-16
C4_102 65 113 7.5e-16
R4_11 64 66 350
C4_111 64 113 1.05e-15
C4_112 66 113 1.05e-15
R4_12 64 79 650
C4_121 64 113 1.95e-15
C4_122 79 113 1.95e-15
R4_13 70 82 700
C4_131 70 113 2.1e-15
C4_132 82 113 2.1e-15
R4_14 58 70 450
C4_141 58 113 1.35e-15
C4_142 70 113 1.35e-15
R4_15 78 79 200
C4_151 78 113 6e-16
C4_152 79 113 6e-16
R4_16 88 92 0.2
C4_161 88 113 7.7e-16
C4_162 92 113 7.7e-16
R4_17 87 88 0.2
C4_171 87 113 7e-16
C4_172 88 113 7e-16
R4_18 76 87 0.5
C4_181 76 113 1.4e-15
C4_182 87 113 1.4e-15
R4_19 63 76 0.5
C4_191 63 113 1.4e-15
C4_192 76 113 1.4e-15
R4_20 81 89 0.6
C4_201 81 113 1.75e-15
C4_202 89 113 1.75e-15
R4_21 69 81 0.4
C4_211 69 113 1.12e-15
C4_212 81 113 1.12e-15
R4_22 59 69 0.5
C4_221 59 113 1.47e-15
C4_222 69 113 1.47e-15
R4_23 80 77 0.1
C4_231 80 113 4.8e-16
C4_232 77 113 4.8e-16
R4_24 68 80 0.05
C4_241 68 113 2.4e-16
C4_242 80 113 2.4e-16
R4_25 71 83 0.2
C4_251 71 113 9.6e-16
C4_252 83 113 9.6e-16
R4_26 67 68 0.85
C4_261 67 113 4.2e-15
C4_262 68 113 4.2e-15
R4_27 71 74 0.35
C4_271 71 113 1.8e-15
C4_272 74 113 1.8e-15
R4_28 75 74 0.05
C4_281 75 113 3.6e-16
C4_282 74 113 3.6e-16
R4_29 67 75 0.05
C4_291 67 113 3.6e-16
C4_292 75 113 3.6e-16
R4_30 91 85 750
C4_301 91 113 2.25e-15
C4_302 85 113 2.25e-15
R4_31 72 90 1
C4_311 72 113 2.87e-15
C4_312 90 113 2.87e-15
R4_32 60 72 0.5
C4_321 60 113 1.47e-15
C4_322 72 113 1.47e-15
R4_33 84 91 450
C4_331 84 113 1.425e-15
C4_332 91 113 1.425e-15
R4_34 73 84 600
C4_341 73 113 1.875e-15
C4_342 84 113 1.875e-15
R4_35 61 73 500
C4_351 61 113 1.5e-15
C4_352 73 113 1.5e-15
R3_1 96 103 0.001
R3_2 95 97 0.001
R3_3 100 101 0.001
C3_31 100 113 3.6e-16
C3_32 101 113 3.6e-16
R3_4 99 100 0.001
C3_41 99 113 7.2e-16
C3_42 100 113 7.2e-16
R3_5 99 107 0.001
C3_51 99 113 4.8e-16
C3_52 107 113 4.8e-16
R3_6 97 107 0.001
C3_61 97 113 1.08e-15
C3_62 107 113 1.08e-15
R3_7 98 97 0.001
C3_71 98 113 9.6e-16
C3_72 97 113 9.6e-16
R3_8 104 106 0.001
C3_81 104 113 6e-16
C3_82 106 113 6e-16
R3_9 105 104 0.001
C3_91 105 113 7.2e-16
C3_92 104 113 7.2e-16
R3_10 103 105 0.1
C3_101 103 113 1.44e-15
C3_102 105 113 1.44e-15
R3_11 102 103 0.001
C3_111 102 113 8.4e-16
C3_112 103 113 8.4e-16
R3_12 101 102 0.001
C3_121 101 113 2.4e-16
C3_122 102 113 2.4e-16
R2_1 110 111 0.001
R2_2 116 117 0.001
R2_3 119 120 0.001
C2_31 119 113 6e-16
C2_32 120 113 6e-16
R2_4 117 119 0.1
C2_41 117 113 2.16e-15
C2_42 119 113 2.16e-15
R2_5 118 117 0.001
C2_51 118 113 8.4e-16
C2_52 117 113 8.4e-16
R2_6 115 118 0.001
C2_61 115 113 2.4e-16
C2_62 118 113 2.4e-16
R2_7 114 115 0.001
C2_71 114 113 3.6e-16
C2_72 115 113 3.6e-16
R2_8 114 113 0.001
C2_81 114 113 1.2e-15
C2_82 113 113 1.2e-15
R2_9 111 113 0.001
C2_91 111 113 1.08e-15
C2_92 113 113 1.08e-15
R2_10 112 111 0.001
C2_101 112 113 9.6e-16
C2_102 111 113 9.6e-16
R1_1 125 126 0.001
R1_2 144 150 0.001
R1_3 133 132 0.001
R1_4 144 148 0.001
R1_5 134 132 0.001
R1_6 143 142 0.001
R1_7 138 137 0.001
R1_8 141 149 0.001
R1_9 123 124 0.001
R1_10 141 142 0.001
R1_11 137 139 0.001
R1_12 153 147 750
C1_121 153 113 2.25e-15
C1_122 147 113 2.25e-15
R1_13 146 153 450
C1_131 146 113 1.425e-15
C1_132 153 113 1.425e-15
R1_14 139 146 600
C1_141 139 113 1.875e-15
C1_142 146 113 1.875e-15
R1_15 130 139 500
C1_151 130 113 1.5e-15
C1_152 139 113 1.5e-15
R1_16 137 154 1
C1_161 137 113 2.87e-15
C1_162 154 113 2.87e-15
R1_17 131 137 0.5
C1_171 131 113 1.47e-15
C1_172 137 113 1.47e-15
R1_18 149 151 0.2
C1_181 149 113 7.7e-16
C1_182 151 113 7.7e-16
R1_19 142 149 0.3
C1_191 142 113 8.4e-16
C1_192 149 113 8.4e-16
R1_20 124 142 0.9
C1_201 124 113 2.66e-15
C1_202 142 113 2.66e-15
R1_21 129 128 250
C1_211 129 113 7.5e-16
C1_212 128 113 7.5e-16
R1_22 140 138 0.05
C1_221 140 113 3.6e-16
C1_222 138 113 3.6e-16
R1_23 127 129 350
C1_231 127 113 1.05e-15
C1_232 129 113 1.05e-15
R1_24 135 140 0.6
C1_241 135 113 3e-15
C1_242 140 113 3e-15
R1_25 143 145 0.35
C1_251 143 113 1.8e-15
C1_252 145 113 1.8e-15
R1_26 127 136 650
C1_261 127 113 1.95e-15
C1_262 136 113 1.95e-15
R1_27 135 134 0.05
C1_271 135 113 3.6e-16
C1_272 134 113 3.6e-16
R1_28 134 145 0.2
C1_281 134 113 9.6e-16
C1_282 145 113 9.6e-16
R1_29 133 136 200
C1_291 133 113 6e-16
C1_292 136 113 6e-16
R1_30 150 152 0.2
C1_301 150 113 7.7e-16
C1_302 152 113 7.7e-16
R1_31 148 150 0.2
C1_311 148 113 7e-16
C1_312 150 113 7e-16
R1_32 132 148 0.5
C1_321 132 113 1.4e-15
C1_322 148 113 1.4e-15
R1_33 126 132 0.5
C1_331 126 113 1.4e-15
C1_332 132 113 1.4e-15
.ends mux

