module LSHIFT2(input [31:0] data, output [31:0] out);
	assign out = data << 2;
endmodule

