module LSHIFT2_26(input [25:0] entrada, output [27:0] saida);
	assign saida = entrada << 2;
endmodule