module decodificador(a, y);
    input [4:0] a;
    output reg [31:0]  y;

    always_comb
        case(a)
            5'b00000:  y  =  32'b00000000000000000000000000000001;
            5'b00001:  y  =  32'b00000000000000000000000000000010;
            5'b00010:  y  =  32'b00000000000000000000000000000100;
            5'b00011:  y  =  32'b00000000000000000000000000001000;
            5'b00100:  y  =  32'b00000000000000000000000000010000;
            5'b00101:  y  =  32'b00000000000000000000000000100000;
            5'b00110:  y  =  32'b00000000000000000000000001000000;
            5'b00111:  y  =  32'b00000000000000000000000010000000;
            5'b01000:  y  =  32'b00000000000000000000000100000000;
            5'b01001:  y  =  32'b00000000000000000000001000000000;
            5'b01010:  y  =  32'b00000000000000000000010000000000;
            5'b01011:  y  =  32'b00000000000000000000100000000000;
            5'b01100:  y  =  32'b00000000000000000001000000000000;
            5'b01101:  y  =  32'b00000000000000000010000000000000;
            5'b01110:  y  =  32'b00000000000000000100000000000000;
            5'b01111:  y  =  32'b00000000000000001000000000000000;
            5'b10000:  y  =  32'b00000000000000010000000000000000;
            5'b10001:  y  =  32'b00000000000000100000000000000000;
            5'b10010:  y  =  32'b00000000000001000000000000000000;
            5'b10011:  y  =  32'b00000000000010000000000000000000;
            5'b10100:  y  =  32'b00000000000100000000000000000000;
            5'b10101:  y  =  32'b00000000001000000000000000000000;
            5'b10110:  y  =  32'b00000000010000000000000000000000;
            5'b10111:  y  =  32'b00000000100000000000000000000000;
            5'b11000:  y  =  32'b00000001000000000000000000000000;
            5'b11001:  y  =  32'b00000010000000000000000000000000;
            5'b11010:  y  =  32'b00000100000000000000000000000000;
            5'b11011:  y  =  32'b00001000000000000000000000000000;
            5'b11100:  y  =  32'b00010000000000000000000000000000;
            5'b11101:  y  =  32'b00100000000000000000000000000000;
            5'b11110:  y  =  32'b01000000000000000000000000000000;
            5'b11111:  y  =  32'b10000000000000000000000000000000;
            default:   y  =  32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
        endcase
endmodule
